library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_program is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_program is
	type rom is array(0 to  24575) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"00",X"32",X"00",X"A0",X"C3",X"66",X"02",X"3A",X"07",X"60",X"0F",X"D0",X"33",X"33",X"C9",
		X"3A",X"00",X"62",X"0F",X"D8",X"33",X"33",X"C9",X"21",X"09",X"60",X"35",X"C8",X"33",X"33",X"C9",
		X"21",X"08",X"60",X"35",X"28",X"F2",X"E1",X"C9",X"87",X"E1",X"5F",X"16",X"00",X"C3",X"32",X"00",
		X"18",X"12",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"11",X"04",X"00",X"06",X"0A",X"79",X"86",X"77",
		X"19",X"10",X"FA",X"C9",X"21",X"27",X"62",X"46",X"0F",X"10",X"FD",X"D8",X"E1",X"C9",X"11",X"08",
		X"69",X"01",X"28",X"00",X"ED",X"B0",X"C9",X"3A",X"18",X"60",X"21",X"1A",X"60",X"86",X"21",X"19",
		X"60",X"86",X"32",X"18",X"60",X"C9",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",
		X"00",X"A0",X"CD",X"5B",X"01",X"E6",X"01",X"C2",X"00",X"40",X"21",X"38",X"01",X"CD",X"6F",X"01",
		X"3A",X"07",X"60",X"A7",X"C2",X"B5",X"00",X"3A",X"26",X"60",X"A7",X"C2",X"98",X"00",X"3A",X"0E",
		X"60",X"A7",X"C2",X"42",X"01",X"00",X"00",X"00",X"CD",X"55",X"01",X"47",X"E6",X"0F",X"4F",X"3A",
		X"11",X"60",X"2F",X"A0",X"E6",X"10",X"17",X"17",X"17",X"B1",X"60",X"6F",X"22",X"10",X"60",X"78",
		X"CB",X"77",X"C2",X"00",X"00",X"21",X"1A",X"60",X"35",X"CD",X"57",X"00",X"CD",X"7B",X"01",X"CD",
		X"E0",X"00",X"21",X"D2",X"00",X"E5",X"3A",X"05",X"60",X"EF",X"C3",X"01",X"3C",X"07",X"B2",X"08",
		X"FE",X"06",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3E",X"01",X"32",X"00",X"A0",X"F1",X"C9",
		X"21",X"80",X"60",X"3A",X"07",X"60",X"A7",X"C0",X"06",X"08",X"16",X"00",X"7E",X"A7",X"28",X"10",
		X"06",X"08",X"21",X"80",X"60",X"36",X"00",X"23",X"10",X"FB",X"7A",X"CD",X"95",X"4A",X"18",X"04",
		X"14",X"2C",X"10",X"E8",X"C3",X"00",X"4A",X"C5",X"CD",X"5B",X"01",X"C1",X"C9",X"7C",X"21",X"88",
		X"60",X"AF",X"BE",X"CA",X"18",X"01",X"35",X"3C",X"32",X"80",X"7D",X"C9",X"06",X"08",X"AF",X"21",
		X"00",X"7D",X"11",X"80",X"60",X"77",X"12",X"2C",X"1C",X"10",X"FA",X"06",X"04",X"12",X"1C",X"10",
		X"FC",X"32",X"80",X"7D",X"32",X"00",X"7C",X"C9",X"53",X"00",X"69",X"80",X"41",X"00",X"70",X"80",
		X"81",X"C9",X"3A",X"00",X"A8",X"CD",X"78",X"3F",X"C3",X"9B",X"00",X"CB",X"10",X"CB",X"10",X"CB",
		X"10",X"E6",X"06",X"02",X"C9",X"3A",X"00",X"A0",X"C3",X"78",X"3F",X"3A",X"00",X"B8",X"2F",X"47",
		X"E6",X"03",X"20",X"04",X"78",X"E6",X"0C",X"C9",X"0E",X"80",X"78",X"E6",X"0C",X"B1",X"C9",X"21",
		X"70",X"69",X"11",X"80",X"98",X"C3",X"00",X"3F",X"ED",X"B0",X"C9",X"CD",X"5B",X"01",X"CB",X"7F",
		X"21",X"03",X"60",X"C2",X"89",X"01",X"36",X"01",X"C9",X"7E",X"A7",X"C8",X"E5",X"3A",X"05",X"60",
		X"FE",X"03",X"CA",X"9D",X"01",X"CD",X"1C",X"01",X"3E",X"03",X"32",X"83",X"60",X"E1",X"36",X"00",
		X"2B",X"34",X"11",X"24",X"60",X"1A",X"96",X"C0",X"77",X"13",X"2B",X"EB",X"1A",X"FE",X"90",X"D0",
		X"86",X"27",X"12",X"11",X"00",X"04",X"CD",X"9F",X"30",X"C9",X"00",X"37",X"00",X"AA",X"AA",X"AA",
		X"50",X"76",X"00",X"CD",X"74",X"08",X"21",X"BA",X"01",X"11",X"B2",X"60",X"01",X"09",X"00",X"ED",
		X"B0",X"3E",X"01",X"32",X"07",X"60",X"32",X"29",X"62",X"32",X"28",X"62",X"CD",X"B8",X"06",X"CD",
		X"07",X"02",X"3E",X"01",X"CD",X"C9",X"49",X"32",X"05",X"60",X"32",X"27",X"62",X"AF",X"32",X"0A",
		X"60",X"CD",X"53",X"0A",X"11",X"04",X"03",X"CD",X"9F",X"30",X"11",X"02",X"02",X"CD",X"9F",X"30",
		X"11",X"00",X"02",X"CD",X"9F",X"30",X"C9",X"3A",X"00",X"B0",X"4F",X"21",X"20",X"60",X"E6",X"03",
		X"C6",X"03",X"77",X"23",X"79",X"0F",X"0F",X"E6",X"03",X"47",X"3E",X"07",X"CA",X"26",X"02",X"3E",
		X"05",X"C6",X"05",X"27",X"10",X"FB",X"77",X"23",X"79",X"01",X"01",X"01",X"11",X"02",X"01",X"E6",
		X"70",X"17",X"17",X"17",X"17",X"CA",X"47",X"02",X"DA",X"41",X"02",X"3C",X"4F",X"5A",X"C3",X"47",
		X"02",X"C6",X"02",X"47",X"57",X"87",X"5F",X"72",X"23",X"73",X"23",X"70",X"23",X"71",X"23",X"3A",
		X"00",X"B0",X"07",X"3E",X"01",X"DA",X"59",X"02",X"3D",X"77",X"21",X"65",X"35",X"11",X"00",X"61",
		X"01",X"AA",X"00",X"ED",X"B0",X"C9",X"C3",X"C8",X"3F",X"00",X"60",X"AF",X"4F",X"77",X"23",X"0D",
		X"20",X"FB",X"10",X"F8",X"06",X"08",X"21",X"00",X"98",X"4F",X"77",X"23",X"0D",X"20",X"FB",X"10",
		X"F8",X"06",X"04",X"3E",X"FD",X"21",X"00",X"90",X"0E",X"00",X"77",X"23",X"0D",X"20",X"FB",X"10",
		X"F7",X"C3",X"1B",X"3F",X"06",X"40",X"3E",X"FF",X"77",X"23",X"10",X"FC",X"3E",X"C0",X"32",X"B0",
		X"60",X"32",X"B1",X"60",X"AF",X"32",X"83",X"7D",X"32",X"86",X"7D",X"32",X"87",X"7D",X"3C",X"31",
		X"F0",X"6B",X"CD",X"C9",X"49",X"CD",X"1C",X"01",X"3E",X"01",X"32",X"00",X"A0",X"26",X"60",X"3A",
		X"B1",X"60",X"6F",X"7E",X"87",X"30",X"1C",X"CD",X"15",X"03",X"CD",X"50",X"03",X"21",X"19",X"60",
		X"34",X"21",X"83",X"63",X"3A",X"1A",X"60",X"BE",X"28",X"E3",X"77",X"CD",X"7F",X"03",X"CD",X"A2",
		X"03",X"18",X"DA",X"E6",X"1F",X"5F",X"16",X"00",X"36",X"FF",X"2C",X"4E",X"36",X"FF",X"2C",X"7D",
		X"FE",X"C0",X"30",X"02",X"3E",X"C0",X"32",X"B1",X"60",X"79",X"21",X"BD",X"02",X"E5",X"21",X"07",
		X"03",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"1C",X"05",X"9B",X"05",X"C6",X"05",X"E9",X"05",X"11",
		X"06",X"2A",X"06",X"B8",X"06",X"3A",X"1A",X"60",X"47",X"E6",X"0F",X"C0",X"CF",X"3A",X"0D",X"60",
		X"CD",X"47",X"03",X"11",X"E0",X"FF",X"CB",X"60",X"28",X"14",X"3E",X"FD",X"77",X"19",X"77",X"19",
		X"77",X"3A",X"0F",X"60",X"A7",X"C8",X"3A",X"0D",X"60",X"EE",X"01",X"CD",X"47",X"03",X"3C",X"77",
		X"19",X"36",X"25",X"19",X"36",X"20",X"C9",X"21",X"40",X"93",X"A7",X"C8",X"21",X"E0",X"90",X"C9",
		X"3A",X"2D",X"62",X"A7",X"C0",X"21",X"B3",X"60",X"3A",X"0D",X"60",X"A7",X"28",X"03",X"21",X"B6",
		X"60",X"7E",X"E6",X"F0",X"47",X"23",X"7E",X"E6",X"0F",X"B0",X"0F",X"0F",X"0F",X"0F",X"21",X"21",
		X"60",X"BE",X"D8",X"3E",X"01",X"32",X"2D",X"62",X"21",X"28",X"62",X"34",X"C3",X"B8",X"06",X"21",
		X"84",X"63",X"7E",X"34",X"A7",X"C0",X"21",X"81",X"63",X"7E",X"47",X"34",X"E6",X"07",X"C0",X"78",
		X"0F",X"0F",X"0F",X"47",X"3A",X"29",X"62",X"80",X"FE",X"05",X"38",X"02",X"3E",X"05",X"32",X"80",
		X"63",X"C9",X"3E",X"03",X"F7",X"D7",X"3A",X"50",X"63",X"0F",X"D8",X"21",X"B8",X"62",X"35",X"C0",
		X"36",X"04",X"3A",X"B9",X"62",X"0F",X"D0",X"21",X"29",X"6A",X"06",X"40",X"DD",X"21",X"A0",X"66",
		X"0F",X"D2",X"E4",X"03",X"DD",X"36",X"09",X"02",X"DD",X"36",X"0A",X"02",X"04",X"04",X"CD",X"F2",
		X"03",X"21",X"BA",X"62",X"35",X"C0",X"3E",X"01",X"32",X"B9",X"62",X"32",X"A0",X"63",X"3E",X"10",
		X"32",X"BA",X"62",X"C9",X"DD",X"36",X"09",X"02",X"DD",X"36",X"0A",X"00",X"CD",X"F2",X"03",X"C3",
		X"DE",X"03",X"70",X"3A",X"19",X"60",X"0F",X"D8",X"04",X"70",X"C9",X"3A",X"27",X"62",X"FE",X"02",
		X"C2",X"13",X"04",X"21",X"08",X"69",X"3A",X"A3",X"63",X"4F",X"FF",X"CD",X"28",X"47",X"D6",X"3B",
		X"32",X"B7",X"63",X"3A",X"91",X"63",X"A7",X"C2",X"26",X"04",X"3A",X"1A",X"60",X"A7",X"C2",X"86",
		X"04",X"3E",X"01",X"32",X"91",X"63",X"21",X"90",X"63",X"34",X"7E",X"FE",X"80",X"CA",X"64",X"04",
		X"3A",X"93",X"63",X"A7",X"C2",X"86",X"04",X"7E",X"47",X"E6",X"1F",X"C2",X"86",X"04",X"21",X"CF",
		X"39",X"CD",X"31",X"47",X"00",X"21",X"F7",X"39",X"00",X"00",X"00",X"3E",X"03",X"32",X"82",X"60",
		X"3A",X"27",X"62",X"0F",X"00",X"78",X"04",X"0F",X"DA",X"86",X"04",X"21",X"0B",X"69",X"0E",X"FC",
		X"FF",X"C3",X"86",X"04",X"AF",X"77",X"23",X"77",X"3A",X"93",X"63",X"A7",X"C2",X"86",X"04",X"21",
		X"5C",X"38",X"00",X"00",X"00",X"C3",X"50",X"04",X"21",X"08",X"69",X"0E",X"44",X"0F",X"D2",X"85",
		X"04",X"3A",X"B7",X"63",X"4F",X"FF",X"3A",X"90",X"63",X"4F",X"11",X"20",X"00",X"3A",X"27",X"62",
		X"FE",X"04",X"CA",X"BE",X"04",X"79",X"A7",X"CA",X"A1",X"04",X"3E",X"EF",X"CB",X"71",X"C2",X"A3",
		X"04",X"3E",X"FA",X"21",X"A4",X"91",X"CD",X"14",X"05",X"3A",X"05",X"69",X"32",X"05",X"69",X"CB",
		X"71",X"C8",X"47",X"79",X"E6",X"07",X"C0",X"78",X"EE",X"03",X"32",X"05",X"69",X"C9",X"3E",X"FD",
		X"21",X"83",X"91",X"CD",X"14",X"05",X"21",X"83",X"91",X"CD",X"14",X"05",X"CB",X"71",X"CA",X"09",
		X"05",X"3A",X"03",X"62",X"FE",X"80",X"D2",X"F1",X"04",X"3E",X"EF",X"21",X"83",X"91",X"CD",X"14",
		X"05",X"3A",X"01",X"69",X"F6",X"80",X"32",X"01",X"69",X"3A",X"05",X"69",X"F6",X"80",X"C3",X"AC",
		X"04",X"3E",X"EF",X"21",X"83",X"91",X"CD",X"14",X"05",X"3A",X"01",X"69",X"E6",X"7F",X"32",X"01",
		X"69",X"3A",X"05",X"69",X"E6",X"7F",X"C3",X"AC",X"04",X"3A",X"03",X"62",X"FE",X"80",X"D2",X"F9",
		X"04",X"C3",X"E1",X"04",X"06",X"03",X"77",X"19",X"3D",X"10",X"FB",X"C9",X"4F",X"CF",X"CD",X"5F",
		X"05",X"79",X"81",X"81",X"4F",X"21",X"29",X"35",X"06",X"00",X"09",X"A7",X"06",X"03",X"1A",X"8E",
		X"27",X"12",X"13",X"23",X"10",X"F8",X"D5",X"1B",X"3A",X"0D",X"60",X"CD",X"6B",X"05",X"D1",X"1B",
		X"21",X"BA",X"60",X"06",X"03",X"1A",X"BE",X"D8",X"C2",X"50",X"05",X"1B",X"2B",X"10",X"F6",X"C9",
		X"CD",X"5F",X"05",X"21",X"B8",X"60",X"1A",X"77",X"13",X"23",X"10",X"FA",X"C3",X"DA",X"05",X"11",
		X"B2",X"60",X"3A",X"0D",X"60",X"A7",X"C8",X"11",X"B5",X"60",X"C9",X"DD",X"21",X"81",X"93",X"A7",
		X"28",X"0A",X"DD",X"21",X"21",X"91",X"18",X"04",X"DD",X"21",X"41",X"92",X"EB",X"11",X"E0",X"FF",
		X"01",X"04",X"03",X"7E",X"0F",X"0F",X"0F",X"0F",X"CD",X"93",X"05",X"7E",X"CD",X"93",X"05",X"2B",
		X"10",X"F1",X"C9",X"E6",X"0F",X"DD",X"77",X"00",X"DD",X"19",X"C9",X"FE",X"03",X"D2",X"BD",X"05",
		X"F5",X"21",X"B2",X"60",X"A7",X"CA",X"AB",X"05",X"21",X"B5",X"60",X"FE",X"02",X"C2",X"B3",X"05",
		X"21",X"B8",X"60",X"AF",X"77",X"23",X"77",X"23",X"77",X"F1",X"C3",X"C6",X"05",X"3D",X"F5",X"CD",
		X"9B",X"05",X"F1",X"C8",X"18",X"F7",X"FE",X"03",X"CA",X"E0",X"05",X"11",X"B4",X"60",X"A7",X"CA",
		X"D5",X"05",X"11",X"B7",X"60",X"FE",X"02",X"C2",X"6B",X"05",X"11",X"BA",X"60",X"C3",X"78",X"05",
		X"3D",X"F5",X"CD",X"C6",X"05",X"F1",X"C8",X"18",X"F7",X"21",X"4B",X"36",X"87",X"F5",X"E6",X"7F",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"5E",X"23",X"56",X"23",X"01",X"E0",X"FF",X"EB",
		X"1A",X"FE",X"3F",X"CA",X"26",X"00",X"77",X"F1",X"30",X"02",X"36",X"10",X"F5",X"13",X"09",X"18",
		X"EF",X"3A",X"07",X"60",X"0F",X"D0",X"3E",X"05",X"CD",X"E9",X"05",X"21",X"01",X"60",X"11",X"E0",
		X"FF",X"DD",X"21",X"BF",X"90",X"06",X"01",X"C3",X"83",X"05",X"A7",X"CA",X"91",X"06",X"3A",X"8C",
		X"63",X"A7",X"C2",X"A8",X"06",X"3A",X"B8",X"63",X"A7",X"C0",X"3A",X"B0",X"62",X"01",X"0A",X"00",
		X"04",X"91",X"C2",X"40",X"06",X"78",X"07",X"07",X"07",X"07",X"32",X"8C",X"63",X"21",X"4A",X"38",
		X"11",X"45",X"90",X"3E",X"06",X"DD",X"21",X"1D",X"00",X"01",X"03",X"00",X"ED",X"B0",X"DD",X"19",
		X"DD",X"E5",X"D1",X"3D",X"C2",X"55",X"06",X"3A",X"8C",X"63",X"4F",X"E6",X"0F",X"47",X"79",X"0F",
		X"0F",X"0F",X"0F",X"E6",X"0F",X"C2",X"89",X"06",X"3E",X"03",X"32",X"8A",X"60",X"3E",X"00",X"32",
		X"86",X"90",X"00",X"00",X"00",X"80",X"47",X"3E",X"FD",X"32",X"C6",X"90",X"78",X"32",X"A6",X"90",
		X"C9",X"3A",X"8C",X"63",X"47",X"E6",X"0F",X"C5",X"CD",X"1C",X"05",X"C1",X"78",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"0F",X"C6",X"0A",X"C3",X"1C",X"05",X"D6",X"01",X"20",X"05",X"21",X"B8",X"63",X"36",
		X"01",X"27",X"32",X"8C",X"63",X"C3",X"6A",X"06",X"4F",X"CF",X"06",X"06",X"11",X"E0",X"FF",X"21",
		X"83",X"93",X"36",X"FD",X"19",X"10",X"FB",X"3A",X"28",X"62",X"91",X"CA",X"D7",X"06",X"47",X"21",
		X"83",X"93",X"36",X"FF",X"19",X"10",X"FB",X"21",X"E3",X"90",X"36",X"1C",X"21",X"C3",X"90",X"36",
		X"34",X"3A",X"29",X"62",X"FE",X"64",X"38",X"05",X"3E",X"63",X"32",X"29",X"62",X"01",X"0A",X"FF",
		X"04",X"91",X"D2",X"F0",X"06",X"81",X"32",X"83",X"90",X"78",X"32",X"A3",X"90",X"C9",X"3A",X"0A",
		X"60",X"EF",X"86",X"09",X"AB",X"09",X"D6",X"09",X"FE",X"09",X"1B",X"0A",X"37",X"0A",X"63",X"0A",
		X"76",X"0A",X"DA",X"0B",X"00",X"00",X"91",X"0C",X"3C",X"12",X"7A",X"19",X"7C",X"12",X"F2",X"12",
		X"44",X"13",X"8F",X"13",X"A1",X"13",X"AA",X"13",X"BB",X"13",X"1E",X"14",X"86",X"14",X"15",X"16",
		X"6B",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"0A",X"60",X"3A",
		X"01",X"60",X"A7",X"C2",X"5C",X"07",X"7E",X"EF",X"79",X"07",X"63",X"07",X"3C",X"12",X"77",X"19",
		X"7C",X"12",X"C3",X"07",X"CB",X"07",X"4B",X"08",X"00",X"00",X"00",X"00",X"36",X"00",X"21",X"05",
		X"60",X"34",X"C9",X"E7",X"AF",X"32",X"92",X"63",X"32",X"A0",X"63",X"3E",X"01",X"32",X"27",X"62",
		X"32",X"29",X"62",X"32",X"28",X"62",X"C3",X"92",X"0C",X"21",X"86",X"7D",X"36",X"00",X"23",X"36",
		X"00",X"11",X"1B",X"03",X"CD",X"9F",X"30",X"1C",X"CD",X"9F",X"30",X"CD",X"65",X"09",X"21",X"09",
		X"60",X"36",X"02",X"23",X"34",X"CD",X"74",X"08",X"CD",X"53",X"0A",X"3A",X"0F",X"60",X"FE",X"01",
		X"CC",X"EE",X"09",X"ED",X"5B",X"22",X"60",X"21",X"6C",X"91",X"CD",X"AD",X"07",X"73",X"23",X"23",
		X"72",X"7A",X"D6",X"0A",X"C2",X"BC",X"07",X"77",X"3C",X"32",X"8E",X"91",X"11",X"01",X"02",X"CD",
		X"40",X"5A",X"C9",X"CD",X"74",X"08",X"21",X"0A",X"60",X"34",X"C9",X"CD",X"BA",X"5A",X"FE",X"00",
		X"C2",X"2D",X"08",X"3E",X"60",X"32",X"8A",X"63",X"0E",X"5F",X"FE",X"00",X"CA",X"3B",X"08",X"C3",
		X"F2",X"07",X"C2",X"94",X"48",X"3A",X"26",X"60",X"A7",X"C2",X"94",X"48",X"C3",X"50",X"42",X"07",
		X"30",X"02",X"3E",X"01",X"CD",X"7A",X"41",X"21",X"00",X"4F",X"3E",X"B0",X"46",X"23",X"5E",X"23",
		X"56",X"12",X"13",X"10",X"FC",X"23",X"7E",X"FE",X"00",X"C2",X"FA",X"07",X"11",X"1E",X"03",X"CD",
		X"9F",X"30",X"13",X"CD",X"9F",X"30",X"21",X"CF",X"39",X"00",X"00",X"00",X"00",X"CD",X"29",X"46",
		X"21",X"08",X"69",X"0E",X"01",X"FF",X"21",X"0B",X"69",X"0E",X"01",X"FF",X"C9",X"3A",X"8B",X"63",
		X"4F",X"3A",X"8A",X"63",X"3D",X"32",X"8A",X"63",X"C3",X"DA",X"07",X"21",X"09",X"60",X"36",X"02",
		X"23",X"34",X"21",X"8A",X"63",X"36",X"00",X"23",X"36",X"00",X"C9",X"E7",X"CD",X"7D",X"55",X"00",
		X"00",X"C9",X"21",X"00",X"90",X"0E",X"04",X"06",X"00",X"3E",X"FD",X"77",X"23",X"10",X"FC",X"0D",
		X"C2",X"57",X"08",X"21",X"00",X"69",X"0E",X"02",X"06",X"C0",X"AF",X"77",X"23",X"10",X"FC",X"0D",
		X"C2",X"68",X"08",X"C9",X"21",X"04",X"90",X"0E",X"20",X"06",X"1C",X"3E",X"FD",X"11",X"04",X"00",
		X"77",X"23",X"10",X"FC",X"19",X"0D",X"C2",X"79",X"08",X"21",X"22",X"91",X"11",X"20",X"00",X"0E",
		X"02",X"3E",X"FD",X"06",X"0E",X"77",X"19",X"10",X"FC",X"21",X"23",X"91",X"0D",X"C2",X"93",X"08",
		X"CD",X"6A",X"48",X"06",X"00",X"3E",X"00",X"77",X"23",X"10",X"FC",X"06",X"80",X"77",X"23",X"10",
		X"FC",X"C9",X"C3",X"67",X"5A",X"EF",X"BA",X"08",X"F8",X"08",X"CD",X"74",X"08",X"AF",X"32",X"07",
		X"60",X"11",X"0C",X"03",X"CD",X"9F",X"30",X"21",X"0A",X"60",X"34",X"CD",X"65",X"09",X"AF",X"C3",
		X"F6",X"56",X"77",X"2C",X"77",X"06",X"04",X"1E",X"09",X"3A",X"01",X"60",X"FE",X"01",X"CA",X"E4",
		X"08",X"06",X"0C",X"1C",X"3A",X"1A",X"60",X"E6",X"07",X"C2",X"F3",X"08",X"7B",X"CD",X"E9",X"05",
		X"CD",X"16",X"06",X"CD",X"07",X"01",X"A0",X"C9",X"CD",X"D5",X"08",X"FE",X"04",X"CA",X"06",X"09",
		X"FE",X"08",X"CA",X"19",X"09",X"C9",X"CD",X"77",X"09",X"21",X"48",X"60",X"06",X"08",X"AF",X"77",
		X"2C",X"10",X"FC",X"21",X"00",X"00",X"C3",X"38",X"09",X"CD",X"77",X"09",X"CD",X"77",X"09",X"11",
		X"48",X"60",X"3A",X"20",X"60",X"12",X"1C",X"21",X"5E",X"09",X"01",X"07",X"00",X"ED",X"B0",X"11",
		X"01",X"01",X"CD",X"9F",X"30",X"21",X"00",X"01",X"22",X"0E",X"60",X"CD",X"74",X"08",X"11",X"40",
		X"60",X"3A",X"20",X"60",X"12",X"1C",X"21",X"5E",X"09",X"01",X"07",X"00",X"ED",X"B0",X"11",X"00",
		X"01",X"CD",X"9F",X"30",X"AF",X"32",X"0A",X"60",X"3E",X"03",X"32",X"05",X"60",X"C9",X"01",X"65",
		X"3A",X"01",X"00",X"00",X"00",X"11",X"00",X"04",X"CD",X"9F",X"30",X"11",X"14",X"03",X"06",X"06",
		X"CD",X"9F",X"30",X"1C",X"10",X"FA",X"C9",X"21",X"01",X"60",X"3E",X"99",X"86",X"27",X"77",X"11",
		X"00",X"04",X"CD",X"9F",X"30",X"C9",X"CD",X"52",X"08",X"CD",X"1C",X"01",X"11",X"82",X"7D",X"CD",
		X"C9",X"49",X"21",X"0A",X"60",X"3A",X"0E",X"60",X"A7",X"C2",X"9F",X"09",X"36",X"01",X"C9",X"3A",
		X"26",X"60",X"3D",X"CA",X"CF",X"48",X"AF",X"CD",X"50",X"48",X"C9",X"21",X"40",X"60",X"11",X"28",
		X"62",X"01",X"08",X"00",X"ED",X"B0",X"2A",X"2A",X"62",X"7E",X"32",X"27",X"62",X"3A",X"0F",X"60",
		X"A7",X"21",X"09",X"60",X"11",X"0A",X"60",X"CA",X"D0",X"09",X"36",X"78",X"EB",X"36",X"02",X"C9",
		X"36",X"01",X"EB",X"36",X"05",X"C9",X"AF",X"32",X"86",X"7D",X"32",X"87",X"7D",X"11",X"02",X"03",
		X"CD",X"9F",X"30",X"11",X"01",X"02",X"CD",X"9F",X"30",X"3E",X"05",X"32",X"0A",X"60",X"3E",X"02",
		X"32",X"E0",X"90",X"3E",X"25",X"32",X"C0",X"90",X"3E",X"20",X"32",X"A0",X"90",X"C9",X"CD",X"EE",
		X"48",X"11",X"28",X"62",X"01",X"08",X"00",X"ED",X"B0",X"2A",X"2A",X"62",X"7E",X"32",X"27",X"62",
		X"3E",X"78",X"32",X"09",X"60",X"3E",X"04",X"32",X"0A",X"60",X"C9",X"AF",X"32",X"86",X"7D",X"32",
		X"87",X"7D",X"11",X"03",X"03",X"CD",X"9F",X"30",X"11",X"01",X"02",X"CD",X"9F",X"30",X"CD",X"EE",
		X"09",X"3E",X"05",X"32",X"0A",X"60",X"C9",X"11",X"04",X"03",X"CD",X"9F",X"30",X"11",X"02",X"02",
		X"CD",X"9F",X"30",X"11",X"00",X"02",X"CD",X"9F",X"30",X"11",X"00",X"06",X"CD",X"9F",X"30",X"21",
		X"0A",X"60",X"34",X"3E",X"01",X"32",X"40",X"93",X"3E",X"25",X"32",X"20",X"93",X"3E",X"20",X"CD",
		X"1F",X"40",X"C9",X"DF",X"CD",X"74",X"08",X"21",X"09",X"60",X"36",X"01",X"2C",X"34",X"11",X"2C",
		X"62",X"1A",X"A7",X"C0",X"34",X"C9",X"3A",X"85",X"63",X"EF",X"8A",X"0A",X"BF",X"0A",X"E8",X"0A",
		X"69",X"30",X"06",X"0B",X"69",X"30",X"68",X"0B",X"B3",X"0B",X"AF",X"32",X"86",X"7D",X"3C",X"32",
		X"87",X"7D",X"11",X"0D",X"38",X"CD",X"A7",X"0D",X"3E",X"FD",X"32",X"A3",X"92",X"32",X"63",X"92",
		X"3E",X"D4",X"32",X"AA",X"91",X"AF",X"32",X"AF",X"62",X"21",X"B4",X"38",X"22",X"C2",X"63",X"21",
		X"CB",X"38",X"22",X"C4",X"63",X"3E",X"40",X"32",X"09",X"60",X"21",X"85",X"63",X"34",X"C9",X"DF",
		X"CD",X"DB",X"4F",X"CD",X"32",X"3F",X"21",X"72",X"69",X"0E",X"30",X"FF",X"21",X"73",X"69",X"0E",
		X"99",X"FF",X"3E",X"1F",X"32",X"8E",X"63",X"AF",X"32",X"76",X"69",X"21",X"8A",X"60",X"36",X"01",
		X"23",X"36",X"03",X"21",X"85",X"63",X"34",X"C9",X"CD",X"6F",X"30",X"3A",X"AF",X"62",X"E6",X"0F",
		X"CC",X"4A",X"30",X"3A",X"73",X"69",X"FE",X"5D",X"D0",X"3E",X"20",X"32",X"09",X"60",X"21",X"85",
		X"63",X"34",X"22",X"C0",X"63",X"C9",X"3A",X"1A",X"60",X"0F",X"D8",X"2A",X"C2",X"63",X"7E",X"FE",
		X"7F",X"CA",X"1E",X"0B",X"23",X"22",X"C2",X"63",X"4F",X"21",X"73",X"69",X"FF",X"C9",X"21",X"5C",
		X"38",X"CD",X"32",X"3F",X"11",X"00",X"69",X"CD",X"00",X"40",X"00",X"00",X"21",X"72",X"69",X"0E",
		X"50",X"FF",X"21",X"73",X"69",X"0E",X"FC",X"FF",X"CD",X"4A",X"30",X"3A",X"8E",X"63",X"FE",X"0A",
		X"C2",X"38",X"0B",X"3E",X"03",X"32",X"82",X"60",X"11",X"2C",X"39",X"CD",X"A7",X"0D",X"3E",X"FD",
		X"32",X"AA",X"90",X"32",X"8A",X"90",X"3E",X"05",X"32",X"8D",X"63",X"3E",X"20",X"32",X"09",X"60",
		X"21",X"85",X"63",X"34",X"22",X"C0",X"63",X"C9",X"3A",X"1A",X"60",X"0F",X"D8",X"2A",X"C4",X"63",
		X"7E",X"FE",X"7F",X"CA",X"86",X"0B",X"23",X"22",X"C4",X"63",X"21",X"73",X"69",X"4F",X"FF",X"21",
		X"72",X"69",X"0E",X"FF",X"FF",X"C9",X"21",X"CB",X"38",X"22",X"C4",X"63",X"3E",X"03",X"32",X"82",
		X"60",X"21",X"DC",X"38",X"3A",X"8D",X"63",X"3D",X"07",X"07",X"07",X"07",X"5F",X"16",X"00",X"19",
		X"EB",X"CD",X"A7",X"0D",X"21",X"8D",X"63",X"35",X"C0",X"3E",X"B0",X"32",X"09",X"60",X"21",X"85",
		X"63",X"34",X"C9",X"21",X"8A",X"60",X"3A",X"09",X"60",X"FE",X"90",X"20",X"0B",X"36",X"0F",X"23",
		X"36",X"03",X"21",X"19",X"81",X"34",X"18",X"09",X"FE",X"18",X"20",X"05",X"21",X"19",X"69",X"35",
		X"00",X"DF",X"AF",X"32",X"85",X"63",X"34",X"23",X"34",X"C9",X"CD",X"1C",X"01",X"DF",X"CD",X"70",
		X"46",X"16",X"06",X"CD",X"F1",X"40",X"5F",X"CD",X"9F",X"30",X"21",X"86",X"7D",X"36",X"01",X"23",
		X"36",X"00",X"21",X"8A",X"60",X"36",X"02",X"23",X"36",X"03",X"21",X"A7",X"63",X"36",X"00",X"21",
		X"DC",X"92",X"22",X"A8",X"63",X"3A",X"2E",X"62",X"FE",X"06",X"38",X"05",X"3E",X"05",X"32",X"2E",
		X"62",X"3A",X"2F",X"62",X"47",X"3A",X"2A",X"62",X"B8",X"28",X"04",X"21",X"2E",X"62",X"34",X"32",
		X"2F",X"62",X"3A",X"2E",X"62",X"47",X"21",X"BC",X"91",X"0E",X"50",X"71",X"0C",X"2B",X"71",X"0C",
		X"2B",X"71",X"0C",X"2B",X"71",X"79",X"FE",X"67",X"CA",X"43",X"0C",X"0C",X"11",X"23",X"00",X"19",
		X"C3",X"2B",X"0C",X"3A",X"A7",X"63",X"3C",X"32",X"A7",X"63",X"3D",X"CB",X"27",X"CB",X"27",X"E5",
		X"CD",X"3D",X"48",X"C5",X"DD",X"2A",X"A8",X"63",X"4F",X"06",X"00",X"09",X"7E",X"DD",X"77",X"60",
		X"23",X"7E",X"DD",X"77",X"40",X"23",X"7E",X"DD",X"77",X"20",X"DD",X"36",X"E0",X"1D",X"C1",X"DD",
		X"E5",X"E1",X"11",X"FC",X"FF",X"19",X"22",X"A8",X"63",X"E1",X"11",X"5F",X"FF",X"19",X"05",X"C2",
		X"29",X"0C",X"11",X"07",X"03",X"CD",X"9F",X"30",X"21",X"09",X"60",X"36",X"A0",X"23",X"34",X"34",
		X"C9",X"DF",X"CD",X"74",X"08",X"AF",X"32",X"8C",X"63",X"11",X"01",X"05",X"CD",X"9F",X"30",X"21",
		X"86",X"7D",X"36",X"00",X"23",X"36",X"01",X"CD",X"20",X"48",X"3D",X"CA",X"D4",X"0C",X"3D",X"CA",
		X"DF",X"0C",X"3D",X"CA",X"F2",X"0C",X"CD",X"43",X"0D",X"21",X"86",X"7D",X"36",X"01",X"3E",X"0B",
		X"32",X"89",X"60",X"11",X"8B",X"3C",X"CD",X"A7",X"0D",X"3A",X"27",X"62",X"FE",X"04",X"CC",X"00",
		X"0D",X"C3",X"A0",X"3F",X"11",X"E4",X"3A",X"3E",X"08",X"32",X"89",X"60",X"C3",X"C6",X"0C",X"11",
		X"5D",X"3B",X"21",X"86",X"7D",X"36",X"01",X"23",X"36",X"00",X"3E",X"09",X"32",X"89",X"60",X"C3",
		X"C6",X"0C",X"CD",X"27",X"0D",X"3E",X"0A",X"32",X"89",X"60",X"11",X"E5",X"3B",X"C3",X"C6",X"0C",
		X"06",X"08",X"21",X"17",X"0D",X"3E",X"FD",X"5E",X"23",X"56",X"23",X"12",X"3E",X"B7",X"13",X"12",
		X"3E",X"FD",X"00",X"00",X"10",X"EF",X"C9",X"CA",X"92",X"CF",X"92",X"D4",X"92",X"D9",X"92",X"2A",
		X"91",X"2F",X"91",X"34",X"91",X"39",X"91",X"21",X"0D",X"93",X"CD",X"30",X"0D",X"21",X"0D",X"92",
		X"06",X"11",X"36",X"FD",X"23",X"10",X"FB",X"CD",X"3E",X"41",X"19",X"06",X"11",X"36",X"68",X"23",
		X"10",X"FB",X"C9",X"21",X"87",X"92",X"CD",X"4C",X"0D",X"21",X"47",X"91",X"06",X"04",X"36",X"FD",
		X"23",X"10",X"FB",X"11",X"1C",X"00",X"19",X"06",X"04",X"36",X"68",X"23",X"10",X"FB",X"C9",X"CD",
		X"56",X"0F",X"CD",X"41",X"24",X"21",X"09",X"60",X"36",X"40",X"23",X"34",X"21",X"5C",X"38",X"00",
		X"00",X"00",X"11",X"00",X"69",X"CD",X"00",X"40",X"00",X"00",X"3A",X"27",X"62",X"FE",X"04",X"28",
		X"0A",X"0F",X"0F",X"D8",X"21",X"0B",X"69",X"0E",X"FC",X"FF",X"C9",X"21",X"08",X"69",X"0E",X"44",
		X"FF",X"11",X"04",X"00",X"01",X"10",X"02",X"21",X"00",X"69",X"CD",X"3D",X"00",X"01",X"F8",X"02",
		X"21",X"03",X"69",X"CD",X"3D",X"00",X"C9",X"1A",X"32",X"B3",X"63",X"FE",X"AA",X"C8",X"13",X"1A",
		X"67",X"44",X"13",X"1A",X"6F",X"4D",X"D5",X"CD",X"F0",X"2F",X"D1",X"22",X"AB",X"63",X"78",X"E6",
		X"07",X"32",X"B4",X"63",X"79",X"E6",X"07",X"32",X"AF",X"63",X"13",X"1A",X"67",X"90",X"D2",X"D3",
		X"0D",X"ED",X"44",X"32",X"B1",X"63",X"13",X"1A",X"6F",X"91",X"32",X"B2",X"63",X"1A",X"E6",X"07",
		X"32",X"B0",X"63",X"D5",X"CD",X"F0",X"2F",X"D1",X"22",X"AD",X"63",X"3A",X"B3",X"63",X"FE",X"02",
		X"F2",X"4F",X"0E",X"3A",X"B2",X"63",X"D6",X"10",X"47",X"3A",X"AF",X"63",X"80",X"32",X"B2",X"63",
		X"3A",X"AF",X"63",X"C6",X"F0",X"2A",X"AB",X"63",X"77",X"2C",X"D6",X"30",X"77",X"3A",X"B3",X"63",
		X"FE",X"01",X"C2",X"19",X"0E",X"AF",X"32",X"B2",X"63",X"3A",X"B2",X"63",X"D6",X"08",X"32",X"B2",
		X"63",X"DA",X"2A",X"0E",X"2C",X"36",X"C0",X"C3",X"19",X"0E",X"3A",X"B0",X"63",X"C6",X"D0",X"2A",
		X"AD",X"63",X"77",X"3A",X"B3",X"63",X"FE",X"01",X"C2",X"3F",X"0E",X"2D",X"36",X"C0",X"2C",X"3A",
		X"B0",X"63",X"FE",X"00",X"CA",X"4B",X"0E",X"C6",X"E0",X"2C",X"77",X"13",X"C3",X"A7",X"0D",X"3A",
		X"B3",X"63",X"FE",X"02",X"C2",X"E8",X"0E",X"3A",X"AF",X"63",X"C6",X"F0",X"32",X"B5",X"63",X"2A",
		X"AB",X"63",X"3A",X"B5",X"63",X"77",X"23",X"7D",X"E6",X"1F",X"CA",X"78",X"0E",X"3A",X"B5",X"63",
		X"FE",X"F0",X"CA",X"78",X"0E",X"D6",X"10",X"77",X"01",X"1F",X"00",X"09",X"3A",X"B1",X"63",X"D6",
		X"08",X"DA",X"CF",X"0E",X"32",X"B1",X"63",X"3A",X"B2",X"63",X"FE",X"00",X"CA",X"62",X"0E",X"3A",
		X"B5",X"63",X"77",X"23",X"7D",X"E6",X"1F",X"CA",X"A0",X"0E",X"3A",X"B5",X"63",X"D6",X"10",X"77",
		X"01",X"1F",X"00",X"09",X"3A",X"B1",X"63",X"D6",X"08",X"DA",X"CF",X"0E",X"32",X"B1",X"63",X"3A",
		X"B2",X"63",X"CB",X"7F",X"C2",X"D3",X"0E",X"3A",X"B5",X"63",X"3C",X"32",X"B5",X"63",X"FE",X"F8",
		X"C2",X"C9",X"0E",X"23",X"3E",X"F0",X"32",X"B5",X"63",X"7D",X"E6",X"1F",X"C2",X"62",X"0E",X"13",
		X"C3",X"A7",X"0D",X"3A",X"B5",X"63",X"3D",X"32",X"B5",X"63",X"FE",X"F0",X"F2",X"E5",X"0E",X"2B",
		X"3E",X"F7",X"32",X"B5",X"63",X"C3",X"62",X"0E",X"3A",X"B3",X"63",X"FE",X"03",X"C2",X"1B",X"0F",
		X"2A",X"AB",X"63",X"3E",X"B3",X"77",X"01",X"20",X"00",X"09",X"3A",X"B1",X"63",X"D6",X"10",X"DA",
		X"14",X"0F",X"32",X"B1",X"63",X"3E",X"B1",X"77",X"01",X"20",X"00",X"09",X"3A",X"B1",X"63",X"D6",
		X"08",X"C3",X"FF",X"0E",X"3E",X"B2",X"77",X"13",X"C3",X"A7",X"0D",X"3A",X"B3",X"63",X"FE",X"07",
		X"F2",X"CF",X"0E",X"FE",X"04",X"CA",X"4C",X"0F",X"FE",X"05",X"CA",X"51",X"0F",X"3E",X"FE",X"32",
		X"B5",X"63",X"2A",X"AB",X"63",X"3A",X"B5",X"63",X"77",X"01",X"20",X"00",X"09",X"3A",X"B1",X"63",
		X"D6",X"08",X"32",X"B1",X"63",X"D2",X"35",X"0F",X"13",X"C3",X"A7",X"0D",X"3E",X"E0",X"C3",X"2F",
		X"0F",X"3E",X"B0",X"C3",X"2F",X"0F",X"06",X"27",X"CD",X"60",X"57",X"AF",X"77",X"2C",X"10",X"FC",
		X"0E",X"0B",X"16",X"80",X"21",X"80",X"62",X"42",X"77",X"23",X"10",X"FC",X"C3",X"E6",X"3F",X"21",
		X"9C",X"3D",X"11",X"80",X"62",X"01",X"40",X"00",X"ED",X"B0",X"3A",X"29",X"62",X"47",X"A7",X"17",
		X"A7",X"17",X"A7",X"17",X"80",X"80",X"C6",X"28",X"FE",X"51",X"38",X"02",X"3E",X"50",X"21",X"B0",
		X"62",X"06",X"03",X"77",X"2C",X"10",X"FC",X"87",X"47",X"3E",X"DC",X"90",X"FE",X"28",X"30",X"02",
		X"3E",X"28",X"77",X"2C",X"77",X"21",X"09",X"62",X"36",X"04",X"2C",X"36",X"08",X"3A",X"27",X"62",
		X"4F",X"CB",X"57",X"20",X"16",X"21",X"00",X"6A",X"3E",X"4F",X"06",X"03",X"77",X"2C",X"36",X"3A",
		X"2C",X"36",X"0F",X"2C",X"36",X"18",X"2C",X"C6",X"10",X"10",X"F1",X"79",X"EF",X"00",X"00",X"D7",
		X"0F",X"1F",X"10",X"87",X"10",X"31",X"11",X"CD",X"00",X"57",X"11",X"A8",X"69",X"CD",X"92",X"40",
		X"00",X"00",X"21",X"EC",X"3D",X"11",X"07",X"64",X"0E",X"1C",X"06",X"05",X"CD",X"2A",X"12",X"21",
		X"F4",X"3D",X"CD",X"FA",X"11",X"21",X"00",X"3E",X"11",X"FC",X"69",X"CD",X"73",X"40",X"00",X"00",
		X"21",X"0C",X"3E",X"CD",X"A6",X"11",X"21",X"1B",X"10",X"11",X"07",X"67",X"01",X"1C",X"08",X"CD",
		X"2A",X"12",X"CD",X"45",X"48",X"06",X"02",X"CD",X"2A",X"12",X"C9",X"00",X"00",X"02",X"02",X"CD",
		X"21",X"47",X"11",X"07",X"64",X"01",X"1C",X"05",X"CD",X"2A",X"12",X"CD",X"86",X"11",X"CD",X"5A",
		X"45",X"11",X"A7",X"65",X"01",X"0C",X"06",X"CD",X"2A",X"12",X"DD",X"21",X"A0",X"65",X"21",X"B8",
		X"69",X"11",X"10",X"00",X"06",X"06",X"CD",X"D3",X"11",X"21",X"FA",X"3D",X"CD",X"FA",X"11",X"21",
		X"04",X"3E",X"11",X"FC",X"69",X"01",X"04",X"00",X"00",X"00",X"21",X"1C",X"3E",X"11",X"44",X"69",
		X"01",X"08",X"00",X"00",X"00",X"21",X"24",X"3E",X"11",X"E4",X"69",X"01",X"18",X"00",X"ED",X"B0",
		X"21",X"10",X"3E",X"CD",X"A6",X"11",X"21",X"3C",X"3E",X"11",X"0C",X"6A",X"01",X"0C",X"00",X"ED",
		X"B0",X"3E",X"01",X"CD",X"D8",X"44",X"C9",X"21",X"EC",X"3D",X"11",X"07",X"64",X"01",X"1C",X"05",
		X"CD",X"2A",X"12",X"CD",X"41",X"47",X"21",X"00",X"66",X"11",X"10",X"00",X"3E",X"01",X"06",X"06",
		X"77",X"19",X"10",X"FC",X"0E",X"02",X"3E",X"08",X"06",X"03",X"21",X"0D",X"66",X"77",X"19",X"10",
		X"FC",X"3E",X"08",X"0D",X"C2",X"A8",X"10",X"21",X"64",X"3E",X"11",X"03",X"66",X"01",X"0E",X"06",
		X"CD",X"EC",X"11",X"21",X"60",X"3E",X"11",X"07",X"66",X"01",X"0C",X"06",X"CD",X"2A",X"12",X"DD",
		X"21",X"00",X"66",X"21",X"84",X"69",X"06",X"06",X"11",X"10",X"00",X"CD",X"D3",X"11",X"21",X"48",
		X"3E",X"11",X"0C",X"6A",X"01",X"0C",X"00",X"ED",X"B0",X"CD",X"DF",X"44",X"00",X"DD",X"36",X"00",
		X"01",X"DD",X"36",X"03",X"58",X"DD",X"36",X"0E",X"58",X"DD",X"36",X"05",X"80",X"DD",X"36",X"0F",
		X"80",X"DD",X"36",X"20",X"01",X"DD",X"36",X"23",X"EB",X"DD",X"36",X"2E",X"EB",X"DD",X"36",X"25",
		X"60",X"DD",X"36",X"2F",X"60",X"11",X"70",X"69",X"21",X"21",X"11",X"01",X"10",X"00",X"00",X"00",
		X"C9",X"37",X"45",X"0F",X"60",X"37",X"45",X"8F",X"F7",X"77",X"45",X"0F",X"60",X"77",X"45",X"8F",
		X"F7",X"CD",X"48",X"47",X"11",X"07",X"64",X"01",X"1C",X"05",X"CD",X"2A",X"12",X"21",X"14",X"3E",
		X"CD",X"A6",X"11",X"21",X"54",X"3E",X"11",X"0C",X"6A",X"01",X"0C",X"00",X"ED",X"B0",X"21",X"82",
		X"11",X"CD",X"E7",X"44",X"01",X"1E",X"02",X"CD",X"EC",X"11",X"21",X"7E",X"11",X"11",X"A7",X"64",
		X"01",X"1C",X"02",X"CD",X"2A",X"12",X"DD",X"21",X"A0",X"64",X"DD",X"36",X"00",X"01",X"DD",X"36",
		X"20",X"01",X"21",X"50",X"69",X"06",X"02",X"11",X"20",X"00",X"CD",X"D3",X"11",X"C9",X"3F",X"0C",
		X"08",X"08",X"73",X"50",X"8D",X"50",X"21",X"A2",X"11",X"11",X"07",X"65",X"01",X"0C",X"0A",X"CD",
		X"2A",X"12",X"DD",X"21",X"00",X"65",X"21",X"7C",X"69",X"06",X"02",X"11",X"10",X"00",X"CD",X"D3",
		X"11",X"C9",X"3B",X"1C",X"02",X"02",X"11",X"83",X"66",X"01",X"0E",X"02",X"CD",X"EC",X"11",X"21",
		X"08",X"3E",X"11",X"87",X"66",X"01",X"0C",X"02",X"CD",X"2A",X"12",X"DD",X"21",X"80",X"66",X"DD",
		X"36",X"00",X"01",X"DD",X"36",X"10",X"01",X"21",X"8C",X"69",X"06",X"02",X"11",X"10",X"00",X"CD",
		X"FA",X"42",X"C9",X"DD",X"7E",X"07",X"77",X"2C",X"DD",X"7E",X"08",X"77",X"2C",X"DD",X"7E",X"03",
		X"77",X"2C",X"DD",X"7E",X"05",X"77",X"2C",X"DD",X"19",X"10",X"E8",X"C9",X"7E",X"12",X"23",X"1C",
		X"1C",X"7E",X"12",X"23",X"7B",X"81",X"5F",X"10",X"F3",X"C9",X"DD",X"21",X"A0",X"66",X"11",X"28",
		X"6A",X"DD",X"36",X"00",X"01",X"7E",X"DD",X"77",X"03",X"12",X"1C",X"23",X"7E",X"DD",X"77",X"07",
		X"12",X"1C",X"23",X"7E",X"DD",X"77",X"08",X"12",X"1C",X"23",X"7E",X"DD",X"77",X"05",X"12",X"23",
		X"7E",X"DD",X"77",X"09",X"23",X"7E",X"DD",X"77",X"0A",X"C9",X"E5",X"C5",X"06",X"04",X"7E",X"12",
		X"23",X"1C",X"10",X"FA",X"C1",X"E1",X"7B",X"81",X"5F",X"10",X"EF",X"C9",X"DF",X"3A",X"27",X"62",
		X"FE",X"03",X"01",X"16",X"E0",X"CA",X"4B",X"12",X"01",X"3F",X"F0",X"DD",X"21",X"00",X"62",X"21",
		X"70",X"69",X"DD",X"36",X"00",X"01",X"DD",X"71",X"03",X"36",X"80",X"2C",X"DD",X"36",X"07",X"80",
		X"36",X"19",X"2C",X"DD",X"36",X"08",X"19",X"71",X"2C",X"DD",X"70",X"05",X"70",X"DD",X"36",X"0F",
		X"01",X"21",X"0A",X"60",X"34",X"11",X"01",X"06",X"CD",X"9F",X"30",X"C9",X"CD",X"BD",X"1D",X"3A",
		X"9D",X"63",X"EF",X"8B",X"12",X"AC",X"12",X"DE",X"12",X"00",X"00",X"DF",X"21",X"70",X"69",X"36",
		X"2A",X"2C",X"36",X"09",X"00",X"21",X"9D",X"63",X"34",X"3E",X"0D",X"32",X"9E",X"63",X"3E",X"08",
		X"32",X"09",X"60",X"CD",X"BD",X"30",X"3E",X"03",X"32",X"88",X"60",X"C9",X"DF",X"3E",X"08",X"32",
		X"09",X"60",X"21",X"9E",X"63",X"35",X"CA",X"CB",X"12",X"21",X"70",X"69",X"7E",X"1F",X"3E",X"02",
		X"1F",X"47",X"AE",X"77",X"2C",X"78",X"E6",X"80",X"AE",X"77",X"C9",X"21",X"70",X"69",X"36",X"2E",
		X"2C",X"36",X"09",X"00",X"21",X"9D",X"63",X"34",X"3E",X"80",X"32",X"09",X"60",X"C9",X"DF",X"CD",
		X"DB",X"30",X"21",X"0A",X"60",X"3A",X"0E",X"60",X"A7",X"CA",X"ED",X"12",X"34",X"34",X"2B",X"36",
		X"01",X"C9",X"CD",X"B8",X"57",X"AF",X"32",X"2C",X"62",X"21",X"28",X"62",X"35",X"7E",X"11",X"40",
		X"60",X"01",X"08",X"00",X"ED",X"B0",X"A7",X"C2",X"34",X"13",X"3E",X"01",X"21",X"B2",X"60",X"CD",
		X"CA",X"13",X"21",X"D4",X"92",X"3A",X"0F",X"60",X"A7",X"28",X"07",X"11",X"02",X"03",X"CD",X"9F",
		X"30",X"2B",X"CD",X"26",X"18",X"11",X"00",X"03",X"CD",X"9F",X"30",X"21",X"09",X"60",X"36",X"C0",
		X"23",X"36",X"10",X"C9",X"0E",X"08",X"3A",X"0F",X"60",X"A7",X"CA",X"3F",X"13",X"0E",X"17",X"79",
		X"32",X"0A",X"60",X"C9",X"CD",X"1C",X"01",X"AF",X"32",X"2C",X"62",X"21",X"28",X"62",X"35",X"7E",
		X"11",X"48",X"60",X"01",X"08",X"00",X"ED",X"B0",X"A7",X"C2",X"7F",X"13",X"3E",X"03",X"21",X"B5",
		X"60",X"CD",X"CA",X"13",X"11",X"03",X"03",X"CD",X"9F",X"30",X"11",X"00",X"03",X"CD",X"9F",X"30",
		X"21",X"D3",X"92",X"CD",X"26",X"18",X"21",X"09",X"60",X"36",X"C0",X"23",X"36",X"11",X"C9",X"0E",
		X"17",X"3A",X"40",X"60",X"A7",X"C2",X"8A",X"13",X"0E",X"08",X"79",X"32",X"0A",X"60",X"C9",X"C3",
		X"85",X"45",X"3A",X"48",X"60",X"34",X"A7",X"C2",X"9C",X"13",X"0E",X"14",X"79",X"32",X"0A",X"60",
		X"C9",X"C3",X"87",X"46",X"3A",X"40",X"60",X"C3",X"4D",X"44",X"3A",X"26",X"60",X"CD",X"60",X"48",
		X"AF",X"32",X"0A",X"60",X"21",X"01",X"01",X"22",X"0D",X"60",X"C9",X"AF",X"32",X"0D",X"60",X"32",
		X"0E",X"60",X"32",X"0A",X"60",X"3C",X"CD",X"F5",X"48",X"C9",X"11",X"C6",X"61",X"12",X"CF",X"13",
		X"01",X"03",X"00",X"ED",X"B0",X"06",X"03",X"21",X"B1",X"61",X"1B",X"1A",X"0F",X"0F",X"0F",X"0F",
		X"E6",X"0F",X"77",X"23",X"1A",X"E6",X"0F",X"77",X"23",X"10",X"EF",X"06",X"0E",X"36",X"10",X"23",
		X"10",X"FB",X"36",X"3F",X"06",X"05",X"21",X"A5",X"61",X"11",X"C7",X"61",X"1A",X"96",X"23",X"13",
		X"1A",X"9E",X"23",X"13",X"1A",X"9E",X"D8",X"C5",X"06",X"19",X"4E",X"1A",X"77",X"79",X"12",X"2B",
		X"1B",X"10",X"F7",X"01",X"F5",X"FF",X"09",X"EB",X"09",X"EB",X"C1",X"10",X"DF",X"C9",X"CD",X"16",
		X"06",X"DF",X"CD",X"74",X"08",X"3E",X"00",X"32",X"0E",X"60",X"32",X"0D",X"60",X"21",X"1C",X"61",
		X"11",X"22",X"00",X"06",X"05",X"3E",X"01",X"BE",X"CA",X"59",X"14",X"19",X"10",X"F9",X"21",X"1C",
		X"61",X"06",X"05",X"3E",X"03",X"BE",X"CA",X"4F",X"14",X"19",X"10",X"F9",X"C3",X"75",X"14",X"3E",
		X"01",X"32",X"0E",X"60",X"32",X"0D",X"60",X"3E",X"00",X"21",X"26",X"60",X"B6",X"CD",X"60",X"48",
		X"3E",X"00",X"32",X"09",X"60",X"21",X"0A",X"60",X"34",X"11",X"0D",X"03",X"06",X"0C",X"CD",X"9F",
		X"30",X"13",X"10",X"FA",X"C9",X"3E",X"01",X"CD",X"C9",X"49",X"32",X"05",X"60",X"32",X"07",X"60",
		X"3E",X"00",X"32",X"0A",X"60",X"C9",X"CD",X"12",X"48",X"21",X"09",X"60",X"7E",X"A7",X"C2",X"DC",
		X"14",X"32",X"86",X"7D",X"32",X"87",X"7D",X"36",X"01",X"21",X"30",X"60",X"36",X"0A",X"23",X"36",
		X"00",X"23",X"36",X"10",X"23",X"36",X"3C",X"23",X"36",X"3E",X"23",X"36",X"00",X"21",X"E8",X"91",
		X"22",X"36",X"60",X"21",X"1C",X"61",X"3A",X"0E",X"60",X"07",X"3C",X"4F",X"11",X"22",X"00",X"06",
		X"04",X"7E",X"B9",X"CA",X"C9",X"14",X"19",X"10",X"F8",X"22",X"38",X"60",X"11",X"F3",X"FF",X"19",
		X"22",X"3A",X"60",X"06",X"00",X"3A",X"35",X"60",X"4F",X"CD",X"FA",X"15",X"21",X"34",X"60",X"35",
		X"C2",X"FC",X"14",X"36",X"3E",X"2B",X"35",X"CA",X"C6",X"15",X"7E",X"06",X"FF",X"04",X"D6",X"0A",
		X"D2",X"ED",X"14",X"C6",X"0A",X"32",X"52",X"91",X"78",X"32",X"72",X"91",X"21",X"30",X"60",X"46",
		X"36",X"0A",X"3A",X"10",X"60",X"CB",X"7F",X"C2",X"46",X"15",X"E6",X"03",X"C2",X"14",X"15",X"3C",
		X"77",X"C3",X"8A",X"15",X"05",X"CA",X"1D",X"15",X"78",X"77",X"C3",X"8A",X"15",X"CB",X"4F",X"C2",
		X"39",X"15",X"3A",X"35",X"60",X"3C",X"FE",X"1E",X"C2",X"2D",X"15",X"3E",X"00",X"32",X"35",X"60",
		X"4F",X"06",X"00",X"CD",X"FA",X"15",X"C3",X"8A",X"15",X"3A",X"35",X"60",X"D6",X"01",X"F2",X"2D",
		X"15",X"3E",X"1D",X"C3",X"2D",X"15",X"3A",X"35",X"60",X"FE",X"1C",X"CA",X"6D",X"15",X"FE",X"1D",
		X"CA",X"C6",X"15",X"2A",X"36",X"60",X"01",X"68",X"90",X"A7",X"ED",X"42",X"CA",X"8A",X"15",X"09",
		X"C6",X"11",X"77",X"01",X"E0",X"FF",X"09",X"22",X"36",X"60",X"C3",X"8A",X"15",X"2A",X"36",X"60",
		X"01",X"20",X"00",X"09",X"A7",X"01",X"08",X"92",X"ED",X"42",X"C2",X"86",X"15",X"21",X"E8",X"91",
		X"3E",X"FD",X"77",X"C3",X"67",X"15",X"09",X"C3",X"80",X"15",X"21",X"32",X"60",X"35",X"C2",X"F9",
		X"15",X"3A",X"31",X"60",X"A7",X"C2",X"B8",X"15",X"3E",X"01",X"32",X"31",X"60",X"11",X"BF",X"01",
		X"FD",X"2A",X"38",X"60",X"FD",X"6E",X"04",X"FD",X"66",X"05",X"E5",X"DD",X"E1",X"CD",X"7C",X"05",
		X"3E",X"10",X"32",X"32",X"60",X"C3",X"F9",X"15",X"AF",X"32",X"31",X"60",X"ED",X"5B",X"38",X"60",
		X"13",X"13",X"13",X"C3",X"A0",X"15",X"ED",X"5B",X"38",X"60",X"AF",X"12",X"21",X"09",X"60",X"36",
		X"80",X"23",X"35",X"06",X"0C",X"21",X"E8",X"91",X"FD",X"2A",X"3A",X"60",X"11",X"E0",X"FF",X"7E",
		X"FD",X"77",X"00",X"FD",X"23",X"19",X"10",X"F7",X"06",X"05",X"11",X"14",X"03",X"CD",X"9F",X"30",
		X"13",X"10",X"FA",X"11",X"1A",X"03",X"CD",X"9F",X"30",X"C9",X"D5",X"E5",X"CB",X"21",X"21",X"0F",
		X"36",X"09",X"EB",X"21",X"74",X"69",X"36",X"24",X"23",X"36",X"0C",X"23",X"1A",X"77",X"13",X"23",
		X"1A",X"77",X"E1",X"D1",X"C9",X"CD",X"BD",X"30",X"3A",X"27",X"62",X"0F",X"D2",X"2F",X"16",X"3A",
		X"88",X"63",X"EF",X"54",X"16",X"70",X"16",X"8A",X"16",X"32",X"17",X"57",X"17",X"8E",X"17",X"0F",
		X"D2",X"41",X"16",X"3A",X"88",X"63",X"EF",X"A3",X"16",X"BB",X"16",X"32",X"17",X"57",X"17",X"8E",
		X"17",X"CD",X"BD",X"1D",X"3A",X"88",X"63",X"EF",X"B6",X"17",X"69",X"30",X"39",X"18",X"6F",X"18",
		X"80",X"18",X"C6",X"18",X"CD",X"08",X"17",X"21",X"5C",X"38",X"CD",X"32",X"3F",X"3E",X"20",X"32",
		X"09",X"60",X"21",X"88",X"63",X"34",X"3E",X"01",X"F7",X"21",X"73",X"69",X"0E",X"FC",X"FF",X"C9",
		X"DF",X"21",X"32",X"39",X"CD",X"32",X"3F",X"3E",X"20",X"32",X"09",X"60",X"21",X"88",X"63",X"34",
		X"3E",X"04",X"F7",X"21",X"73",X"69",X"0E",X"04",X"FF",X"C9",X"DF",X"21",X"8C",X"38",X"CD",X"32",
		X"3F",X"3E",X"66",X"32",X"76",X"69",X"AF",X"32",X"8E",X"69",X"00",X"00",X"00",X"32",X"AF",X"62",
		X"C3",X"62",X"16",X"CD",X"08",X"17",X"3A",X"7A",X"69",X"D6",X"3B",X"21",X"5C",X"38",X"CD",X"32",
		X"3F",X"21",X"72",X"69",X"4F",X"FF",X"21",X"88",X"63",X"34",X"C9",X"AF",X"32",X"A0",X"62",X"3A",
		X"A3",X"63",X"4F",X"3A",X"7A",X"69",X"FE",X"5A",X"D2",X"E1",X"16",X"CB",X"79",X"CA",X"D5",X"16",
		X"3E",X"01",X"32",X"A0",X"62",X"CD",X"02",X"26",X"3A",X"A3",X"63",X"4F",X"21",X"72",X"69",X"FF",
		X"C9",X"FE",X"5D",X"DA",X"EE",X"16",X"CB",X"79",X"CA",X"D0",X"16",X"C3",X"D5",X"16",X"21",X"8C",
		X"38",X"CD",X"32",X"3F",X"3E",X"66",X"32",X"76",X"69",X"AF",X"32",X"8E",X"69",X"00",X"00",X"00",
		X"32",X"AF",X"62",X"21",X"88",X"63",X"34",X"C9",X"CD",X"1C",X"01",X"C3",X"13",X"17",X"36",X"80",
		X"23",X"36",X"76",X"CD",X"F0",X"45",X"CD",X"35",X"40",X"21",X"05",X"69",X"36",X"10",X"21",X"83",
		X"91",X"11",X"20",X"00",X"3E",X"FD",X"CD",X"14",X"05",X"21",X"8A",X"60",X"36",X"07",X"23",X"36",
		X"03",X"C9",X"CD",X"A0",X"59",X"3A",X"7B",X"69",X"FE",X"2C",X"D0",X"CD",X"0A",X"41",X"AF",X"32",
		X"04",X"69",X"32",X"76",X"69",X"3E",X"6B",X"32",X"8E",X"69",X"3D",X"00",X"00",X"00",X"CD",X"54",
		X"40",X"00",X"21",X"88",X"63",X"34",X"C9",X"CD",X"6F",X"30",X"CD",X"E1",X"45",X"00",X"00",X"CD",
		X"83",X"17",X"3E",X"40",X"32",X"09",X"60",X"21",X"88",X"63",X"34",X"C9",X"11",X"03",X"00",X"21",
		X"8F",X"69",X"06",X"08",X"C3",X"CC",X"45",X"52",X"FE",X"19",X"D2",X"7F",X"17",X"36",X"00",X"2B",
		X"10",X"F2",X"C9",X"06",X"08",X"7E",X"A7",X"C2",X"26",X"00",X"19",X"10",X"F8",X"C9",X"DF",X"2A",
		X"2A",X"62",X"23",X"7E",X"FE",X"7F",X"C2",X"9D",X"17",X"21",X"75",X"3A",X"7E",X"22",X"2A",X"62",
		X"32",X"27",X"62",X"11",X"00",X"05",X"CD",X"9F",X"30",X"AF",X"32",X"88",X"63",X"21",X"09",X"60",
		X"36",X"30",X"23",X"36",X"08",X"C9",X"00",X"CD",X"1C",X"01",X"21",X"8A",X"60",X"36",X"0E",X"23",
		X"36",X"03",X"3E",X"FD",X"11",X"20",X"00",X"21",X"23",X"92",X"00",X"00",X"00",X"21",X"83",X"91",
		X"CD",X"14",X"05",X"21",X"DA",X"92",X"CD",X"26",X"18",X"11",X"47",X"3A",X"CD",X"A7",X"0D",X"21",
		X"D5",X"92",X"CD",X"26",X"18",X"11",X"4D",X"3A",X"CD",X"A7",X"0D",X"21",X"D0",X"92",X"CD",X"26",
		X"18",X"11",X"53",X"3A",X"CD",X"A7",X"0D",X"21",X"CB",X"92",X"CD",X"26",X"18",X"11",X"59",X"3A",
		X"CD",X"A7",X"0D",X"21",X"5C",X"38",X"CD",X"32",X"48",X"21",X"72",X"69",X"0E",X"44",X"FF",X"21",
		X"05",X"69",X"36",X"13",X"3E",X"20",X"32",X"09",X"60",X"3E",X"80",X"32",X"90",X"63",X"21",X"88",
		X"63",X"34",X"22",X"C0",X"63",X"C9",X"11",X"DB",X"FF",X"0E",X"0E",X"3E",X"10",X"06",X"05",X"77",
		X"23",X"10",X"FC",X"19",X"0D",X"C2",X"2D",X"18",X"C9",X"CD",X"65",X"41",X"34",X"CA",X"59",X"18",
		X"7E",X"E6",X"07",X"C0",X"11",X"CF",X"39",X"CB",X"5E",X"20",X"03",X"11",X"F7",X"39",X"EB",X"CD",
		X"32",X"3F",X"21",X"72",X"69",X"0E",X"44",X"FF",X"C9",X"21",X"5C",X"38",X"CD",X"32",X"3F",X"21",
		X"72",X"69",X"0E",X"44",X"FF",X"98",X"99",X"32",X"09",X"60",X"21",X"88",X"63",X"34",X"C9",X"DF",
		X"21",X"1F",X"3A",X"CD",X"32",X"3F",X"9B",X"03",X"32",X"84",X"60",X"21",X"88",X"63",X"34",X"C9",
		X"21",X"73",X"69",X"0E",X"01",X"FF",X"3A",X"83",X"69",X"FE",X"D0",X"C0",X"3E",X"20",X"32",X"80",
		X"69",X"21",X"24",X"6A",X"36",X"7F",X"2C",X"36",X"39",X"2C",X"36",X"01",X"2C",X"36",X"D8",X"21",
		X"C6",X"92",X"CD",X"26",X"18",X"11",X"5F",X"3A",X"CD",X"A7",X"0D",X"11",X"04",X"00",X"01",X"28",
		X"02",X"21",X"03",X"69",X"CD",X"3D",X"00",X"3E",X"00",X"32",X"AF",X"62",X"3E",X"03",X"32",X"82",
		X"60",X"CD",X"C0",X"57",X"34",X"C9",X"CD",X"05",X"19",X"35",X"CA",X"3D",X"19",X"7E",X"E6",X"07",
		X"C0",X"CD",X"44",X"44",X"7E",X"EE",X"80",X"77",X"21",X"19",X"69",X"46",X"CB",X"A8",X"AF",X"CD",
		X"09",X"30",X"F6",X"20",X"77",X"21",X"AF",X"62",X"7E",X"FE",X"E0",X"C2",X"10",X"19",X"3E",X"50",
		X"32",X"8B",X"69",X"C3",X"70",X"55",X"FF",X"FF",X"3E",X"9F",X"32",X"8A",X"69",X"3A",X"03",X"62",
		X"FE",X"80",X"C3",X"0F",X"19",X"CD",X"0C",X"40",X"21",X"AF",X"62",X"C9",X"32",X"8A",X"69",X"7E",
		X"FE",X"C0",X"C0",X"21",X"8A",X"60",X"36",X"0C",X"3A",X"29",X"62",X"0F",X"38",X"02",X"36",X"05",
		X"23",X"36",X"03",X"21",X"23",X"6A",X"36",X"40",X"2B",X"36",X"09",X"2B",X"36",X"76",X"2B",X"36",
		X"8F",X"3A",X"03",X"62",X"FE",X"80",X"D0",X"3E",X"6F",X"32",X"20",X"6A",X"C9",X"2A",X"2A",X"62",
		X"23",X"7E",X"FE",X"7F",X"C2",X"4B",X"19",X"21",X"75",X"3A",X"7E",X"22",X"2A",X"62",X"32",X"27",
		X"62",X"21",X"29",X"62",X"34",X"11",X"00",X"05",X"CD",X"9F",X"30",X"AF",X"32",X"2E",X"62",X"32",
		X"88",X"63",X"21",X"09",X"60",X"36",X"E0",X"23",X"36",X"08",X"C9",X"CD",X"52",X"08",X"3A",X"0E",
		X"60",X"C6",X"12",X"32",X"0A",X"60",X"C9",X"CD",X"EE",X"21",X"CD",X"BD",X"1D",X"CD",X"8C",X"1E",
		X"CD",X"C3",X"1A",X"CD",X"72",X"1F",X"CD",X"8F",X"2C",X"CD",X"03",X"2C",X"CD",X"ED",X"30",X"CD",
		X"04",X"2E",X"CD",X"EA",X"24",X"CD",X"DB",X"2D",X"CD",X"D4",X"2E",X"CD",X"07",X"22",X"CD",X"33",
		X"1A",X"CD",X"85",X"2A",X"CD",X"46",X"1F",X"CD",X"FA",X"26",X"CD",X"F2",X"25",X"CD",X"DA",X"19",
		X"CD",X"FB",X"03",X"CD",X"08",X"28",X"CD",X"1D",X"28",X"CD",X"57",X"1E",X"CD",X"07",X"1A",X"CD",
		X"CB",X"2F",X"00",X"00",X"00",X"3A",X"00",X"62",X"A7",X"C0",X"CD",X"1C",X"01",X"21",X"82",X"60",
		X"36",X"03",X"21",X"0A",X"60",X"34",X"2B",X"36",X"40",X"C9",X"3A",X"03",X"62",X"06",X"03",X"21",
		X"0C",X"6A",X"BE",X"CA",X"ED",X"19",X"2C",X"2C",X"2C",X"2C",X"10",X"F6",X"C9",X"3A",X"05",X"62",
		X"2C",X"2C",X"2C",X"BE",X"C0",X"2D",X"2D",X"CB",X"5E",X"C0",X"2D",X"CD",X"EE",X"44",X"AF",X"32",
		X"42",X"63",X"3C",X"32",X"40",X"63",X"C9",X"3A",X"86",X"63",X"EF",X"1E",X"1A",X"15",X"1A",X"1F",
		X"1A",X"2A",X"1A",X"00",X"00",X"AF",X"32",X"87",X"63",X"3E",X"02",X"32",X"86",X"63",X"C9",X"21",
		X"87",X"63",X"35",X"C0",X"3E",X"03",X"32",X"86",X"63",X"C9",X"3A",X"16",X"62",X"A7",X"C0",X"E1",
		X"C3",X"D2",X"19",X"3E",X"08",X"F7",X"3A",X"03",X"62",X"FE",X"4B",X"CA",X"4B",X"1A",X"FE",X"B3",
		X"CA",X"4B",X"1A",X"3A",X"91",X"62",X"3D",X"CA",X"51",X"1A",X"C9",X"3E",X"01",X"32",X"91",X"62",
		X"C9",X"32",X"91",X"62",X"47",X"3A",X"05",X"62",X"3D",X"FE",X"D0",X"D0",X"07",X"D2",X"62",X"1A",
		X"CB",X"D0",X"07",X"07",X"D2",X"69",X"1A",X"CB",X"C8",X"E6",X"07",X"FE",X"06",X"C2",X"72",X"1A",
		X"CB",X"C8",X"3A",X"03",X"62",X"07",X"D2",X"7B",X"1A",X"CB",X"C0",X"21",X"92",X"62",X"78",X"85",
		X"6F",X"7E",X"A7",X"C8",X"36",X"00",X"21",X"90",X"62",X"35",X"78",X"01",X"05",X"00",X"1F",X"DA",
		X"BD",X"1A",X"21",X"CB",X"02",X"A7",X"CA",X"9E",X"1A",X"09",X"3D",X"C2",X"99",X"1A",X"01",X"00",
		X"90",X"09",X"3E",X"10",X"77",X"2D",X"77",X"2C",X"2C",X"77",X"3E",X"01",X"32",X"40",X"63",X"32",
		X"42",X"63",X"32",X"25",X"62",X"3A",X"16",X"62",X"A7",X"CC",X"95",X"1D",X"C9",X"21",X"2B",X"01",
		X"C3",X"95",X"1A",X"3A",X"16",X"62",X"3D",X"CA",X"B2",X"1B",X"3A",X"1E",X"62",X"A7",X"C2",X"55",
		X"1B",X"3A",X"17",X"62",X"3D",X"CA",X"E6",X"1A",X"3A",X"15",X"62",X"3D",X"CA",X"38",X"1B",X"3A",
		X"10",X"60",X"17",X"DA",X"6E",X"1B",X"CD",X"1F",X"24",X"3A",X"10",X"60",X"1D",X"CA",X"F5",X"1A",
		X"CB",X"47",X"C2",X"8F",X"1C",X"15",X"CA",X"FE",X"1A",X"CB",X"4F",X"C2",X"AB",X"1C",X"3A",X"17",
		X"62",X"3D",X"C8",X"3A",X"05",X"62",X"C6",X"08",X"57",X"3A",X"03",X"62",X"F6",X"03",X"CB",X"97",
		X"01",X"15",X"00",X"CD",X"6E",X"23",X"F5",X"21",X"07",X"62",X"7E",X"E6",X"80",X"F6",X"06",X"77",
		X"21",X"1A",X"62",X"3E",X"04",X"B9",X"36",X"01",X"D2",X"2C",X"1B",X"35",X"F1",X"A7",X"CA",X"4E",
		X"1B",X"7E",X"A7",X"C0",X"2C",X"72",X"2C",X"70",X"3A",X"10",X"60",X"CB",X"5F",X"C2",X"F2",X"1C",
		X"3A",X"15",X"62",X"A7",X"C8",X"3A",X"10",X"60",X"CB",X"57",X"C2",X"03",X"1D",X"C9",X"2C",X"70",
		X"2C",X"72",X"C3",X"45",X"1B",X"21",X"1E",X"62",X"35",X"C0",X"3A",X"18",X"62",X"32",X"17",X"62",
		X"21",X"07",X"62",X"7E",X"E6",X"80",X"77",X"AF",X"32",X"02",X"62",X"C3",X"A6",X"1D",X"3E",X"01",
		X"32",X"16",X"62",X"21",X"10",X"62",X"3A",X"10",X"60",X"01",X"80",X"00",X"1F",X"DA",X"8A",X"1B",
		X"01",X"80",X"FF",X"1F",X"DA",X"8A",X"1B",X"01",X"00",X"00",X"AF",X"70",X"2C",X"71",X"2C",X"36",
		X"01",X"2C",X"36",X"48",X"2C",X"77",X"32",X"04",X"62",X"32",X"06",X"62",X"3A",X"07",X"62",X"E6",
		X"80",X"F6",X"0E",X"32",X"07",X"62",X"3A",X"05",X"62",X"32",X"0E",X"62",X"21",X"81",X"60",X"36",
		X"03",X"C9",X"DD",X"21",X"00",X"62",X"3A",X"03",X"62",X"DD",X"77",X"0B",X"3A",X"05",X"62",X"DD",
		X"77",X"0C",X"CD",X"9C",X"23",X"CD",X"1F",X"24",X"15",X"C2",X"F2",X"1B",X"DD",X"36",X"10",X"00",
		X"DD",X"36",X"11",X"80",X"DD",X"CB",X"07",X"FE",X"3A",X"20",X"62",X"3D",X"CA",X"EC",X"1B",X"CD",
		X"07",X"24",X"DD",X"74",X"12",X"DD",X"75",X"13",X"DD",X"36",X"14",X"00",X"CD",X"9C",X"23",X"C3",
		X"A6",X"1D",X"1D",X"C2",X"05",X"1C",X"DD",X"36",X"10",X"FF",X"DD",X"36",X"11",X"80",X"DD",X"CB",
		X"07",X"BE",X"C3",X"D8",X"1B",X"CD",X"1C",X"2B",X"3D",X"CA",X"3A",X"1C",X"3A",X"1F",X"62",X"3D",
		X"CA",X"76",X"1C",X"3A",X"14",X"62",X"D6",X"14",X"C2",X"33",X"1C",X"3E",X"01",X"32",X"1F",X"62",
		X"CD",X"53",X"28",X"A7",X"CA",X"A6",X"1D",X"32",X"42",X"63",X"3E",X"01",X"32",X"40",X"63",X"32",
		X"25",X"62",X"00",X"3C",X"CC",X"54",X"29",X"C3",X"A6",X"1D",X"05",X"CA",X"4F",X"1C",X"3C",X"32",
		X"1F",X"62",X"AF",X"21",X"10",X"62",X"06",X"05",X"77",X"2C",X"10",X"FC",X"C3",X"A6",X"1D",X"32",
		X"16",X"62",X"3A",X"20",X"62",X"EE",X"01",X"32",X"00",X"62",X"21",X"07",X"62",X"7E",X"E6",X"80",
		X"F6",X"0F",X"77",X"3E",X"04",X"32",X"1E",X"62",X"AF",X"32",X"1F",X"62",X"3A",X"25",X"62",X"3D",
		X"CC",X"95",X"1D",X"C3",X"A6",X"1D",X"3A",X"05",X"62",X"21",X"0E",X"62",X"D6",X"0F",X"BE",X"DA",
		X"A6",X"1D",X"3E",X"01",X"32",X"20",X"62",X"21",X"84",X"60",X"36",X"03",X"C3",X"A6",X"1D",X"06",
		X"01",X"3A",X"0F",X"62",X"A7",X"C2",X"D2",X"1C",X"3A",X"02",X"62",X"47",X"3E",X"05",X"CD",X"09",
		X"30",X"32",X"02",X"62",X"E6",X"03",X"F6",X"80",X"C3",X"C2",X"1C",X"06",X"FF",X"3A",X"0F",X"62",
		X"A7",X"C2",X"D2",X"1C",X"3A",X"02",X"62",X"47",X"3E",X"01",X"CD",X"09",X"30",X"32",X"02",X"62",
		X"E6",X"03",X"21",X"07",X"62",X"77",X"1F",X"DC",X"8F",X"1D",X"3E",X"02",X"32",X"0F",X"62",X"C3",
		X"A6",X"1D",X"21",X"03",X"62",X"7E",X"80",X"77",X"3A",X"27",X"62",X"3D",X"C2",X"EB",X"1C",X"66",
		X"3A",X"05",X"62",X"6F",X"CD",X"33",X"23",X"7D",X"32",X"05",X"62",X"21",X"0F",X"62",X"35",X"C3",
		X"A6",X"1D",X"3A",X"0F",X"62",X"A7",X"C2",X"8A",X"1D",X"3E",X"03",X"32",X"0F",X"62",X"3E",X"02",
		X"C3",X"11",X"1D",X"3A",X"0F",X"62",X"A7",X"C2",X"76",X"1D",X"3E",X"04",X"32",X"0F",X"62",X"3E",
		X"FE",X"21",X"05",X"62",X"86",X"77",X"47",X"3A",X"22",X"62",X"EE",X"01",X"32",X"22",X"62",X"C2",
		X"51",X"1D",X"78",X"C6",X"08",X"21",X"1C",X"62",X"BE",X"CA",X"67",X"1D",X"2D",X"96",X"CA",X"67",
		X"1D",X"06",X"05",X"D6",X"08",X"CA",X"3F",X"1D",X"05",X"D6",X"04",X"CA",X"3F",X"1D",X"05",X"3E",
		X"80",X"21",X"07",X"62",X"A6",X"EE",X"80",X"B0",X"77",X"3E",X"01",X"32",X"15",X"62",X"C3",X"A6",
		X"1D",X"2D",X"2D",X"7E",X"F6",X"03",X"CB",X"97",X"77",X"3A",X"24",X"62",X"EE",X"01",X"32",X"24",
		X"62",X"CC",X"8F",X"1D",X"C3",X"49",X"1D",X"3E",X"06",X"32",X"07",X"62",X"AF",X"32",X"19",X"62",
		X"32",X"15",X"62",X"C3",X"A6",X"1D",X"3A",X"1A",X"62",X"A7",X"CA",X"8A",X"1D",X"32",X"19",X"62",
		X"3A",X"1C",X"62",X"D6",X"13",X"21",X"05",X"62",X"BE",X"D0",X"21",X"0F",X"62",X"35",X"C9",X"3E",
		X"03",X"32",X"80",X"60",X"C9",X"32",X"25",X"62",X"3A",X"27",X"62",X"3D",X"00",X"21",X"8A",X"60",
		X"36",X"0D",X"2C",X"36",X"03",X"C9",X"21",X"70",X"69",X"3A",X"07",X"62",X"77",X"3A",X"08",X"62",
		X"2C",X"77",X"3A",X"03",X"62",X"2C",X"77",X"3A",X"05",X"62",X"C3",X"80",X"57",X"3A",X"40",X"63",
		X"EF",X"49",X"1E",X"C9",X"1D",X"4A",X"1E",X"00",X"00",X"3E",X"40",X"32",X"41",X"63",X"3E",X"02",
		X"32",X"40",X"63",X"3A",X"42",X"63",X"1F",X"DA",X"70",X"3E",X"1F",X"DA",X"00",X"1E",X"1F",X"DA",
		X"F5",X"1D",X"21",X"85",X"60",X"36",X"03",X"3A",X"29",X"62",X"3D",X"CA",X"00",X"1E",X"3D",X"CA",
		X"08",X"1E",X"C3",X"10",X"1E",X"3A",X"18",X"60",X"1F",X"DA",X"08",X"1E",X"1F",X"DA",X"10",X"1E",
		X"06",X"33",X"11",X"03",X"00",X"C3",X"15",X"1E",X"06",X"36",X"11",X"05",X"00",X"C3",X"15",X"1E",
		X"06",X"37",X"11",X"08",X"00",X"CD",X"9F",X"30",X"2A",X"43",X"63",X"7E",X"36",X"00",X"2C",X"2C",
		X"2C",X"4E",X"C3",X"36",X"1E",X"11",X"01",X"00",X"CD",X"9F",X"30",X"3A",X"05",X"62",X"C6",X"14",
		X"4F",X"3A",X"03",X"62",X"00",X"00",X"21",X"74",X"69",X"70",X"2C",X"36",X"04",X"2C",X"77",X"2C",
		X"71",X"3E",X"05",X"F7",X"21",X"85",X"60",X"36",X"03",X"C9",X"21",X"41",X"63",X"35",X"C0",X"AF",
		X"32",X"76",X"69",X"32",X"40",X"63",X"C9",X"3A",X"27",X"62",X"CB",X"57",X"C2",X"80",X"1E",X"1F",
		X"3A",X"05",X"62",X"DA",X"7A",X"1E",X"FE",X"51",X"D0",X"3A",X"03",X"62",X"17",X"3E",X"00",X"DA",
		X"74",X"1E",X"3E",X"80",X"32",X"70",X"69",X"C3",X"85",X"1E",X"FE",X"31",X"D0",X"C3",X"6D",X"1E",
		X"3A",X"90",X"62",X"A7",X"C0",X"3E",X"16",X"32",X"0A",X"60",X"E1",X"C9",X"3A",X"50",X"63",X"A7",
		X"C8",X"CD",X"96",X"1E",X"E1",X"C9",X"3A",X"45",X"63",X"EF",X"A0",X"1E",X"09",X"1F",X"23",X"1F",
		X"3A",X"52",X"63",X"FE",X"65",X"21",X"80",X"69",X"CA",X"85",X"47",X"21",X"78",X"69",X"DA",X"B4",
		X"1E",X"21",X"7C",X"69",X"DD",X"2A",X"51",X"63",X"16",X"00",X"3A",X"53",X"63",X"5F",X"01",X"04",
		X"00",X"3A",X"54",X"63",X"A7",X"CA",X"CF",X"1E",X"09",X"DD",X"19",X"3D",X"C2",X"C8",X"1E",X"DD",
		X"36",X"00",X"00",X"DD",X"7E",X"15",X"A7",X"3E",X"02",X"CA",X"DE",X"1E",X"3E",X"04",X"32",X"42",
		X"63",X"CD",X"46",X"3F",X"00",X"00",X"00",X"02",X"0C",X"2C",X"3E",X"60",X"02",X"0C",X"2C",X"3E",
		X"0C",X"02",X"0C",X"2C",X"7E",X"02",X"21",X"45",X"63",X"34",X"2C",X"36",X"06",X"2C",X"36",X"05",
		X"21",X"8A",X"60",X"36",X"06",X"2C",X"36",X"03",X"C9",X"21",X"46",X"63",X"35",X"C0",X"36",X"06",
		X"2C",X"35",X"CA",X"1D",X"1F",X"21",X"2D",X"6A",X"7E",X"EE",X"01",X"77",X"C9",X"36",X"04",X"2D",
		X"2D",X"34",X"C9",X"21",X"46",X"63",X"35",X"C0",X"36",X"0C",X"2C",X"35",X"CA",X"34",X"1F",X"21",
		X"2D",X"6A",X"34",X"C9",X"2D",X"2D",X"AF",X"77",X"32",X"50",X"63",X"3C",X"32",X"40",X"63",X"21",
		X"2C",X"6A",X"22",X"43",X"63",X"C9",X"3A",X"21",X"62",X"A7",X"C8",X"AF",X"32",X"04",X"62",X"32",
		X"06",X"62",X"32",X"21",X"62",X"32",X"10",X"62",X"32",X"11",X"62",X"32",X"12",X"62",X"32",X"13",
		X"62",X"32",X"14",X"62",X"3C",X"32",X"16",X"62",X"32",X"1F",X"62",X"3A",X"05",X"62",X"32",X"0E",
		X"62",X"C9",X"3A",X"27",X"62",X"3D",X"C0",X"DD",X"21",X"00",X"67",X"21",X"7C",X"69",X"11",X"20",
		X"00",X"06",X"04",X"DD",X"7E",X"00",X"3D",X"CA",X"93",X"1F",X"2C",X"2C",X"2C",X"2C",X"DD",X"19",
		X"10",X"F1",X"C9",X"DD",X"7E",X"01",X"3D",X"CA",X"EC",X"20",X"DD",X"7E",X"02",X"1F",X"DA",X"AC",
		X"1F",X"1F",X"DA",X"E5",X"1F",X"1F",X"DA",X"EF",X"1F",X"C3",X"53",X"20",X"D9",X"DD",X"34",X"05",
		X"DD",X"7E",X"17",X"DD",X"BE",X"05",X"C2",X"CE",X"1F",X"DD",X"7E",X"15",X"07",X"07",X"C6",X"15",
		X"DD",X"77",X"07",X"DD",X"7E",X"02",X"EE",X"07",X"DD",X"77",X"02",X"C3",X"BA",X"21",X"DD",X"7E",
		X"0F",X"3D",X"C2",X"DF",X"1F",X"DD",X"7E",X"07",X"EE",X"01",X"DD",X"77",X"07",X"3E",X"04",X"DD",
		X"77",X"0F",X"C3",X"BA",X"21",X"D9",X"01",X"00",X"01",X"DD",X"34",X"03",X"C3",X"F6",X"1F",X"D9",
		X"01",X"04",X"FF",X"DD",X"35",X"03",X"DD",X"66",X"03",X"DD",X"6E",X"05",X"7C",X"E6",X"07",X"FE",
		X"03",X"CA",X"5F",X"21",X"2D",X"2D",X"2D",X"CD",X"33",X"23",X"2C",X"2C",X"2C",X"7D",X"DD",X"77",
		X"05",X"CD",X"DE",X"23",X"CD",X"B4",X"24",X"DD",X"7E",X"03",X"FE",X"2A",X"DA",X"2F",X"20",X"FE",
		X"D4",X"DA",X"BA",X"21",X"AF",X"DD",X"77",X"10",X"DD",X"36",X"11",X"60",X"C3",X"38",X"20",X"AF",
		X"DD",X"36",X"10",X"FF",X"DD",X"36",X"11",X"A0",X"DD",X"36",X"12",X"FF",X"DD",X"36",X"13",X"F0",
		X"DD",X"77",X"14",X"DD",X"77",X"0E",X"DD",X"77",X"04",X"DD",X"77",X"06",X"DD",X"36",X"02",X"08",
		X"C3",X"BA",X"21",X"D9",X"CD",X"9C",X"23",X"CD",X"2F",X"2A",X"A7",X"C2",X"83",X"20",X"DD",X"7E",
		X"03",X"C6",X"08",X"FE",X"10",X"DA",X"79",X"20",X"CD",X"B4",X"24",X"DD",X"7E",X"10",X"E6",X"01",
		X"07",X"07",X"4F",X"CD",X"DE",X"23",X"C3",X"BA",X"21",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"03",
		X"C3",X"BA",X"21",X"DD",X"34",X"0E",X"DD",X"7E",X"0E",X"3D",X"CA",X"A2",X"20",X"3D",X"CA",X"C3",
		X"20",X"DD",X"7E",X"10",X"3D",X"3E",X"04",X"C2",X"9C",X"20",X"3E",X"02",X"DD",X"77",X"02",X"C3",
		X"BA",X"21",X"DD",X"7E",X"15",X"A7",X"C2",X"B5",X"20",X"21",X"05",X"62",X"DD",X"7E",X"05",X"D6",
		X"16",X"BE",X"D2",X"C3",X"20",X"DD",X"7E",X"10",X"A7",X"C2",X"E1",X"20",X"DD",X"77",X"11",X"DD",
		X"36",X"10",X"FF",X"CD",X"07",X"24",X"CB",X"3C",X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"DD",X"74",
		X"12",X"DD",X"75",X"13",X"AF",X"DD",X"77",X"14",X"DD",X"77",X"04",X"DD",X"77",X"06",X"C3",X"BA",
		X"21",X"DD",X"36",X"10",X"01",X"DD",X"36",X"11",X"00",X"C3",X"C3",X"20",X"D9",X"CD",X"9C",X"23",
		X"7C",X"D6",X"1A",X"DD",X"46",X"19",X"B8",X"DA",X"04",X"21",X"CD",X"2F",X"2A",X"A7",X"C2",X"18",
		X"21",X"CD",X"B4",X"24",X"DD",X"7E",X"03",X"C6",X"08",X"FE",X"10",X"D2",X"CE",X"1F",X"AF",X"DD",
		X"77",X"00",X"DD",X"77",X"03",X"C3",X"BA",X"21",X"DD",X"7E",X"05",X"FE",X"E0",X"DA",X"46",X"21",
		X"DD",X"7E",X"07",X"E6",X"FC",X"F6",X"01",X"DD",X"77",X"07",X"AF",X"DD",X"77",X"01",X"DD",X"77",
		X"02",X"DD",X"36",X"10",X"FF",X"DD",X"77",X"11",X"DD",X"77",X"12",X"DD",X"36",X"13",X"B0",X"DD",
		X"36",X"0E",X"01",X"C3",X"53",X"21",X"CD",X"07",X"24",X"CD",X"CB",X"22",X"DD",X"7E",X"05",X"DD",
		X"77",X"19",X"AF",X"DD",X"77",X"14",X"DD",X"77",X"04",X"DD",X"77",X"06",X"C3",X"BA",X"21",X"7D",
		X"C6",X"05",X"57",X"7C",X"01",X"15",X"00",X"CD",X"6D",X"21",X"C3",X"BA",X"21",X"CD",X"6E",X"23",
		X"3D",X"C0",X"78",X"D6",X"05",X"DD",X"77",X"17",X"3A",X"48",X"63",X"A7",X"CA",X"B2",X"21",X"3A",
		X"05",X"62",X"D6",X"10",X"BA",X"D8",X"3A",X"80",X"63",X"1F",X"3C",X"47",X"3A",X"18",X"60",X"4F",
		X"E6",X"03",X"B8",X"D0",X"21",X"10",X"60",X"3A",X"03",X"62",X"BB",X"CA",X"B2",X"21",X"D2",X"A9",
		X"21",X"CB",X"46",X"CA",X"AE",X"21",X"C3",X"B2",X"21",X"CB",X"4E",X"C2",X"B2",X"21",X"79",X"E6",
		X"18",X"C0",X"DD",X"34",X"07",X"DD",X"CB",X"02",X"C6",X"C9",X"D9",X"DD",X"7E",X"07",X"77",X"2C",
		X"DD",X"7E",X"08",X"77",X"2C",X"DD",X"7E",X"03",X"77",X"2C",X"DD",X"7E",X"05",X"77",X"C3",X"8D",
		X"1F",X"80",X"FE",X"01",X"3A",X"04",X"30",X"02",X"10",X"82",X"28",X"02",X"10",X"82",X"78",X"01",
		X"10",X"81",X"FF",X"02",X"38",X"01",X"80",X"02",X"FF",X"04",X"80",X"04",X"60",X"80",X"11",X"D1",
		X"21",X"21",X"CC",X"63",X"7E",X"07",X"83",X"5F",X"1A",X"32",X"10",X"60",X"2C",X"7E",X"35",X"A7",
		X"C0",X"1C",X"1A",X"77",X"2D",X"34",X"C9",X"3E",X"02",X"F7",X"3A",X"1A",X"60",X"1F",X"21",X"80",
		X"62",X"7E",X"DA",X"19",X"22",X"21",X"88",X"62",X"7E",X"E5",X"EF",X"27",X"22",X"59",X"22",X"99",
		X"22",X"A2",X"22",X"00",X"00",X"00",X"00",X"E1",X"2C",X"35",X"C2",X"3A",X"22",X"2D",X"34",X"2C",
		X"2C",X"CD",X"43",X"22",X"3E",X"01",X"32",X"1A",X"62",X"C9",X"2C",X"CD",X"43",X"22",X"AF",X"32",
		X"1A",X"62",X"C9",X"3A",X"05",X"62",X"FE",X"7A",X"D2",X"57",X"22",X"3A",X"16",X"62",X"A7",X"C2",
		X"57",X"22",X"3A",X"03",X"62",X"BE",X"C8",X"E1",X"C9",X"E1",X"2C",X"2C",X"2C",X"2C",X"35",X"C0",
		X"3E",X"04",X"77",X"2D",X"34",X"CD",X"BD",X"22",X"3E",X"78",X"BE",X"C2",X"75",X"22",X"2D",X"2D",
		X"2D",X"34",X"2C",X"2C",X"2C",X"2D",X"CD",X"43",X"22",X"3A",X"05",X"62",X"FE",X"68",X"D2",X"8A",
		X"22",X"21",X"05",X"62",X"34",X"CD",X"C0",X"3F",X"34",X"C9",X"1F",X"DA",X"81",X"22",X"1F",X"3E",
		X"01",X"DA",X"95",X"22",X"AF",X"32",X"22",X"62",X"C9",X"E1",X"3A",X"18",X"60",X"E6",X"3C",X"C0",
		X"34",X"C9",X"E1",X"2C",X"2C",X"2C",X"2C",X"35",X"C0",X"36",X"02",X"2D",X"35",X"CD",X"BD",X"22",
		X"3E",X"68",X"BE",X"C0",X"AF",X"06",X"80",X"2D",X"2D",X"70",X"2D",X"77",X"C9",X"7E",X"CB",X"5D",
		X"C3",X"49",X"43",X"C2",X"C9",X"22",X"11",X"47",X"69",X"12",X"C9",X"3A",X"48",X"63",X"A7",X"CA",
		X"E1",X"22",X"3A",X"80",X"63",X"3D",X"EF",X"F6",X"22",X"F6",X"22",X"03",X"23",X"03",X"23",X"1A",
		X"23",X"3A",X"29",X"62",X"47",X"05",X"3E",X"01",X"CA",X"F9",X"22",X"05",X"3E",X"B1",X"CA",X"F9",
		X"22",X"3E",X"E9",X"C3",X"F9",X"22",X"3A",X"18",X"60",X"DD",X"77",X"11",X"E6",X"01",X"3D",X"DD",
		X"77",X"10",X"C9",X"3A",X"18",X"60",X"DD",X"77",X"11",X"3A",X"03",X"62",X"DD",X"BE",X"03",X"3E",
		X"01",X"D2",X"16",X"23",X"3D",X"3D",X"DD",X"77",X"10",X"C9",X"3A",X"03",X"62",X"DD",X"96",X"03",
		X"0E",X"FF",X"DA",X"26",X"23",X"0C",X"07",X"CB",X"11",X"07",X"CB",X"11",X"DD",X"71",X"10",X"DD",
		X"77",X"11",X"C9",X"3E",X"0F",X"A4",X"05",X"CA",X"42",X"23",X"FE",X"0F",X"D8",X"06",X"FF",X"C3",
		X"47",X"23",X"FE",X"01",X"D0",X"06",X"01",X"3E",X"F0",X"BD",X"CA",X"60",X"23",X"3E",X"4C",X"BD",
		X"CA",X"66",X"23",X"7D",X"CB",X"6F",X"CA",X"5C",X"23",X"90",X"6F",X"C9",X"80",X"C3",X"5A",X"23",
		X"CB",X"7C",X"C2",X"59",X"23",X"C9",X"7C",X"FE",X"98",X"D8",X"7D",X"C3",X"5C",X"23",X"21",X"00",
		X"63",X"ED",X"B1",X"C2",X"9A",X"23",X"E5",X"C5",X"01",X"14",X"00",X"09",X"0C",X"5F",X"7A",X"BE",
		X"CA",X"8F",X"23",X"09",X"BE",X"CA",X"95",X"23",X"57",X"7B",X"C1",X"E1",X"C3",X"71",X"23",X"09",
		X"3E",X"01",X"C3",X"98",X"23",X"AF",X"ED",X"42",X"C1",X"46",X"E1",X"C9",X"DD",X"7E",X"04",X"DD",
		X"86",X"11",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"DD",X"8E",X"10",X"DD",X"77",X"03",X"DD",X"7E",
		X"06",X"DD",X"96",X"13",X"6F",X"DD",X"7E",X"05",X"DD",X"9E",X"12",X"67",X"DD",X"7E",X"14",X"A7",
		X"17",X"3C",X"06",X"00",X"CB",X"10",X"CB",X"27",X"CB",X"10",X"CB",X"27",X"CB",X"10",X"CB",X"27",
		X"CB",X"10",X"4F",X"09",X"DD",X"74",X"05",X"DD",X"75",X"06",X"DD",X"34",X"14",X"C9",X"DD",X"7E",
		X"0F",X"3D",X"C2",X"03",X"24",X"AF",X"DD",X"CB",X"07",X"26",X"17",X"DD",X"CB",X"08",X"26",X"17",
		X"47",X"3E",X"03",X"B1",X"CD",X"09",X"30",X"1F",X"DD",X"CB",X"08",X"1E",X"1F",X"DD",X"CB",X"07",
		X"1E",X"3E",X"04",X"DD",X"77",X"0F",X"C9",X"DD",X"7E",X"14",X"07",X"07",X"07",X"07",X"4F",X"E6",
		X"0F",X"67",X"79",X"E6",X"F0",X"6F",X"DD",X"4E",X"13",X"DD",X"46",X"12",X"ED",X"42",X"C9",X"11",
		X"00",X"01",X"3A",X"03",X"62",X"FE",X"16",X"D8",X"15",X"1C",X"FE",X"EA",X"D0",X"1D",X"3A",X"27",
		X"62",X"0F",X"D0",X"3A",X"05",X"62",X"FE",X"58",X"D0",X"3A",X"03",X"62",X"FE",X"6C",X"D0",X"14",
		X"C9",X"21",X"FA",X"37",X"3E",X"5E",X"06",X"06",X"86",X"23",X"10",X"FC",X"FD",X"21",X"10",X"63",
		X"A7",X"CA",X"56",X"24",X"FD",X"23",X"3A",X"27",X"62",X"3D",X"21",X"E4",X"3A",X"CA",X"71",X"24",
		X"3D",X"21",X"5D",X"3B",X"CA",X"71",X"24",X"3D",X"21",X"E5",X"3B",X"CA",X"71",X"24",X"21",X"8B",
		X"3C",X"DD",X"21",X"00",X"63",X"11",X"05",X"00",X"7E",X"A7",X"CA",X"88",X"24",X"3D",X"CA",X"9E",
		X"24",X"FE",X"A9",X"C8",X"19",X"C3",X"78",X"24",X"23",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",
		X"77",X"15",X"23",X"23",X"7E",X"DD",X"77",X"2A",X"DD",X"23",X"23",X"C3",X"78",X"24",X"23",X"7E",
		X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"15",X"23",X"23",X"7E",X"FD",X"77",X"2A",X"FD",X"23",
		X"23",X"C3",X"78",X"24",X"DD",X"7E",X"05",X"FE",X"E8",X"D8",X"DD",X"7E",X"03",X"FE",X"2A",X"D0",
		X"FE",X"20",X"D8",X"DD",X"7E",X"15",X"A7",X"CA",X"D0",X"24",X"3E",X"03",X"32",X"B9",X"62",X"AF",
		X"DD",X"77",X"00",X"DD",X"77",X"03",X"21",X"82",X"60",X"36",X"03",X"E1",X"3A",X"48",X"63",X"A7",
		X"C2",X"BA",X"21",X"3C",X"32",X"48",X"63",X"C3",X"BA",X"21",X"3E",X"02",X"F7",X"CD",X"23",X"25",
		X"CD",X"91",X"25",X"DD",X"21",X"A0",X"65",X"06",X"03",X"21",X"80",X"69",X"DD",X"7E",X"00",X"A7",
		X"CA",X"1C",X"25",X"DD",X"7E",X"07",X"77",X"2C",X"DD",X"7E",X"08",X"77",X"2C",X"DD",X"7E",X"03",
		X"77",X"2C",X"DD",X"7E",X"05",X"77",X"2C",X"DD",X"19",X"10",X"E1",X"C9",X"7D",X"C6",X"04",X"6F",
		X"C3",X"17",X"25",X"21",X"9B",X"63",X"7E",X"A7",X"C2",X"8F",X"25",X"3A",X"9A",X"63",X"A7",X"C8",
		X"06",X"03",X"11",X"10",X"00",X"DD",X"21",X"A0",X"65",X"DD",X"CB",X"00",X"46",X"CA",X"45",X"25",
		X"DD",X"19",X"10",X"F5",X"C9",X"CD",X"57",X"00",X"FE",X"60",X"DD",X"36",X"05",X"7C",X"DA",X"58",
		X"25",X"3A",X"A3",X"62",X"3D",X"C2",X"6E",X"25",X"DD",X"36",X"05",X"CC",X"3A",X"A6",X"62",X"07",
		X"DD",X"36",X"03",X"07",X"D2",X"76",X"25",X"DD",X"36",X"03",X"F8",X"C3",X"76",X"25",X"CD",X"57",
		X"00",X"FE",X"68",X"C3",X"60",X"25",X"DD",X"36",X"00",X"01",X"DD",X"36",X"07",X"3A",X"DD",X"36",
		X"09",X"08",X"DD",X"36",X"0A",X"03",X"3E",X"7C",X"32",X"9B",X"63",X"AF",X"32",X"9A",X"63",X"35",
		X"C9",X"DD",X"21",X"A0",X"65",X"11",X"10",X"00",X"06",X"03",X"DD",X"CB",X"00",X"46",X"CA",X"BB",
		X"25",X"DD",X"7E",X"03",X"67",X"C6",X"07",X"FE",X"0E",X"DA",X"D6",X"25",X"DD",X"7E",X"05",X"FE",
		X"7C",X"CA",X"C0",X"25",X"3A",X"A6",X"63",X"84",X"DD",X"77",X"03",X"DD",X"19",X"10",X"DB",X"C9",
		X"7C",X"FE",X"80",X"CA",X"D6",X"25",X"3A",X"A5",X"63",X"D2",X"CF",X"25",X"3A",X"A4",X"63",X"84",
		X"DD",X"77",X"03",X"C3",X"BB",X"25",X"21",X"80",X"69",X"C3",X"EE",X"42",X"CA",X"E7",X"25",X"2C",
		X"2C",X"2C",X"2C",X"3D",X"C3",X"DC",X"25",X"AF",X"DD",X"77",X"00",X"DD",X"77",X"03",X"00",X"C3",
		X"7D",X"45",X"3E",X"02",X"F7",X"CD",X"02",X"26",X"CD",X"2F",X"26",X"CD",X"79",X"26",X"CD",X"D3",
		X"2A",X"C9",X"3A",X"1A",X"60",X"0F",X"DA",X"16",X"26",X"21",X"A0",X"62",X"35",X"C2",X"16",X"26",
		X"36",X"80",X"2C",X"CD",X"DE",X"26",X"21",X"A1",X"62",X"CD",X"E9",X"26",X"32",X"A3",X"63",X"3A",
		X"1A",X"60",X"E6",X"1F",X"FE",X"01",X"C0",X"11",X"AA",X"93",X"EB",X"CD",X"A6",X"26",X"C9",X"21",
		X"A3",X"62",X"3A",X"05",X"62",X"FE",X"C0",X"DA",X"6F",X"26",X"3A",X"1A",X"60",X"0F",X"DA",X"4C",
		X"26",X"2D",X"35",X"C2",X"4C",X"26",X"36",X"C0",X"2C",X"CD",X"DE",X"26",X"21",X"A3",X"62",X"CD",
		X"E9",X"26",X"32",X"A5",X"63",X"ED",X"44",X"32",X"A4",X"63",X"3A",X"1A",X"60",X"E6",X"1F",X"C0",
		X"2D",X"11",X"CF",X"91",X"EB",X"CD",X"A6",X"26",X"E6",X"7F",X"21",X"ED",X"69",X"77",X"C9",X"CB",
		X"7E",X"C2",X"4C",X"26",X"36",X"FF",X"C3",X"4C",X"26",X"3A",X"1A",X"60",X"0F",X"DA",X"8D",X"26",
		X"21",X"A5",X"62",X"35",X"C2",X"8D",X"26",X"36",X"FF",X"2C",X"CD",X"DE",X"26",X"21",X"A6",X"62",
		X"CD",X"E9",X"26",X"32",X"A6",X"63",X"3A",X"1A",X"60",X"E6",X"1F",X"FE",X"02",X"C0",X"11",X"B9",
		X"93",X"EB",X"CD",X"A6",X"26",X"C9",X"CD",X"2C",X"45",X"DA",X"C5",X"26",X"7E",X"3C",X"FE",X"23",
		X"C2",X"B5",X"26",X"3E",X"20",X"77",X"7D",X"CD",X"44",X"45",X"7E",X"3D",X"FE",X"1F",X"C2",X"C3",
		X"26",X"3E",X"22",X"77",X"C9",X"7E",X"3D",X"FE",X"1F",X"C2",X"CE",X"26",X"3E",X"22",X"77",X"7D",
		X"CD",X"44",X"45",X"7E",X"3C",X"FE",X"23",X"C2",X"DC",X"26",X"3E",X"20",X"77",X"C9",X"CB",X"7E",
		X"CA",X"E6",X"26",X"36",X"02",X"C9",X"36",X"FE",X"C9",X"3A",X"1A",X"60",X"E6",X"01",X"C8",X"C3",
		X"40",X"57",X"FF",X"C2",X"F8",X"26",X"3E",X"01",X"77",X"C9",X"3E",X"04",X"F7",X"3A",X"05",X"62",
		X"FE",X"F0",X"D2",X"7F",X"27",X"3A",X"29",X"62",X"3D",X"3A",X"1A",X"60",X"C2",X"1A",X"27",X"E6",
		X"03",X"FE",X"01",X"CA",X"1E",X"27",X"DA",X"22",X"27",X"C9",X"0F",X"DA",X"22",X"27",X"CD",X"45",
		X"27",X"C9",X"CD",X"97",X"27",X"CD",X"DA",X"27",X"06",X"03",X"11",X"10",X"00",X"21",X"84",X"69",
		X"DD",X"21",X"00",X"66",X"DD",X"7E",X"03",X"2C",X"2C",X"77",X"2C",X"DD",X"7E",X"05",X"77",X"2C",
		X"DD",X"19",X"10",X"F0",X"C9",X"3A",X"98",X"63",X"A7",X"C8",X"3A",X"16",X"62",X"A7",X"C0",X"3A",
		X"03",X"62",X"FE",X"2C",X"DA",X"66",X"27",X"FE",X"43",X"DA",X"6F",X"27",X"FE",X"6C",X"DA",X"66",
		X"27",X"FE",X"83",X"DA",X"87",X"27",X"AF",X"32",X"98",X"63",X"3C",X"32",X"21",X"62",X"C9",X"3A",
		X"05",X"62",X"FE",X"71",X"DA",X"7F",X"27",X"3D",X"32",X"05",X"62",X"32",X"73",X"69",X"C9",X"AF",
		X"32",X"00",X"62",X"32",X"98",X"63",X"C9",X"3A",X"05",X"62",X"FE",X"E8",X"D2",X"7F",X"27",X"3C",
		X"32",X"05",X"62",X"32",X"73",X"69",X"C9",X"06",X"06",X"11",X"10",X"00",X"DD",X"21",X"00",X"66",
		X"DD",X"CB",X"00",X"46",X"CA",X"C2",X"27",X"DD",X"CB",X"0D",X"5E",X"CA",X"C7",X"27",X"DD",X"7E",
		X"05",X"3D",X"DD",X"77",X"05",X"FE",X"60",X"C2",X"C2",X"27",X"DD",X"36",X"03",X"77",X"DD",X"36",
		X"0D",X"04",X"DD",X"19",X"10",X"DA",X"C9",X"DD",X"7E",X"05",X"3C",X"DD",X"77",X"05",X"FE",X"F8",
		X"C2",X"C2",X"27",X"DD",X"36",X"00",X"00",X"C3",X"C2",X"27",X"21",X"A7",X"62",X"7E",X"A7",X"C2",
		X"06",X"28",X"06",X"03",X"DD",X"21",X"00",X"66",X"DD",X"CB",X"00",X"46",X"CA",X"F4",X"27",X"DD",
		X"19",X"10",X"F5",X"C9",X"DD",X"36",X"00",X"01",X"DD",X"36",X"03",X"37",X"DD",X"36",X"05",X"F8",
		X"DD",X"36",X"0D",X"08",X"36",X"34",X"35",X"C9",X"FD",X"21",X"00",X"62",X"3A",X"05",X"62",X"4F",
		X"21",X"07",X"04",X"CD",X"6F",X"28",X"A7",X"C8",X"3D",X"32",X"00",X"62",X"C9",X"06",X"02",X"11",
		X"10",X"00",X"FD",X"21",X"80",X"66",X"FD",X"CB",X"01",X"46",X"C2",X"32",X"28",X"FD",X"19",X"10",
		X"F5",X"C9",X"FD",X"4E",X"05",X"FD",X"66",X"09",X"FD",X"6E",X"0A",X"CD",X"6F",X"28",X"A7",X"C8",
		X"32",X"50",X"63",X"3A",X"B9",X"63",X"90",X"32",X"54",X"63",X"7B",X"32",X"53",X"63",X"DD",X"22",
		X"51",X"63",X"C9",X"FD",X"21",X"00",X"62",X"3A",X"05",X"62",X"C6",X"0C",X"4F",X"3A",X"10",X"60",
		X"E6",X"03",X"21",X"08",X"05",X"CA",X"6B",X"28",X"21",X"08",X"13",X"CD",X"88",X"3E",X"C9",X"3A",
		X"27",X"62",X"E5",X"EF",X"00",X"00",X"80",X"28",X"B0",X"28",X"E0",X"28",X"01",X"29",X"00",X"00",
		X"E1",X"06",X"04",X"78",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"67",X"CD",X"13",
		X"29",X"CD",X"E9",X"42",X"32",X"B9",X"63",X"1E",X"20",X"DD",X"21",X"00",X"64",X"CD",X"13",X"29",
		X"06",X"01",X"78",X"32",X"B9",X"63",X"1E",X"00",X"DD",X"21",X"A0",X"66",X"CD",X"13",X"29",X"C9",
		X"E1",X"CD",X"E9",X"42",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"64",X"CD",X"13",
		X"29",X"06",X"03",X"78",X"32",X"B9",X"63",X"1E",X"10",X"DD",X"21",X"A0",X"65",X"CD",X"13",X"29",
		X"06",X"01",X"78",X"32",X"B9",X"63",X"1E",X"00",X"DD",X"21",X"A0",X"66",X"CD",X"13",X"29",X"C9",
		X"E1",X"CD",X"E9",X"42",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"64",X"CD",X"13",
		X"29",X"06",X"0A",X"78",X"32",X"B9",X"63",X"1E",X"10",X"DD",X"21",X"00",X"65",X"CD",X"13",X"29",
		X"C9",X"E1",X"CD",X"E9",X"42",X"32",X"B9",X"63",X"11",X"20",X"00",X"DD",X"21",X"00",X"64",X"CD",
		X"13",X"29",X"C9",X"DD",X"E5",X"DD",X"CB",X"00",X"46",X"CA",X"4C",X"29",X"79",X"DD",X"96",X"05",
		X"D2",X"25",X"29",X"ED",X"44",X"3C",X"95",X"DA",X"30",X"29",X"DD",X"96",X"0A",X"D2",X"4C",X"29",
		X"FD",X"7E",X"03",X"DD",X"96",X"03",X"D2",X"3B",X"29",X"ED",X"44",X"94",X"DA",X"45",X"29",X"DD",
		X"96",X"09",X"D2",X"4C",X"29",X"3E",X"01",X"DD",X"E1",X"33",X"33",X"C9",X"DD",X"19",X"10",X"C5",
		X"AF",X"DD",X"E1",X"C9",X"3E",X"0B",X"F7",X"CD",X"74",X"29",X"32",X"18",X"62",X"0F",X"0F",X"32",
		X"85",X"60",X"78",X"A7",X"C8",X"FE",X"01",X"CA",X"6F",X"29",X"DD",X"36",X"01",X"01",X"C9",X"DD",
		X"36",X"11",X"01",X"C9",X"FD",X"21",X"00",X"62",X"3A",X"05",X"62",X"4F",X"21",X"08",X"04",X"06",
		X"02",X"11",X"10",X"00",X"DD",X"21",X"80",X"66",X"CD",X"13",X"29",X"C9",X"2A",X"C8",X"63",X"7D",
		X"C6",X"0E",X"6F",X"56",X"2C",X"7E",X"C6",X"0C",X"5F",X"EB",X"CD",X"F0",X"2F",X"7E",X"FE",X"B0",
		X"DA",X"AC",X"29",X"E6",X"0F",X"FE",X"08",X"D2",X"AC",X"29",X"AF",X"C9",X"3E",X"01",X"C9",X"3E",
		X"04",X"F7",X"FD",X"21",X"00",X"62",X"3A",X"05",X"62",X"4F",X"21",X"08",X"04",X"CD",X"22",X"2A",
		X"A7",X"CA",X"20",X"2A",X"3E",X"06",X"90",X"CA",X"D0",X"29",X"DD",X"19",X"3D",X"C3",X"C7",X"29",
		X"DD",X"7E",X"05",X"D6",X"04",X"57",X"3A",X"0C",X"62",X"C6",X"05",X"BA",X"D2",X"EE",X"29",X"7A",
		X"D6",X"08",X"32",X"05",X"62",X"3E",X"01",X"47",X"32",X"98",X"63",X"33",X"33",X"C9",X"3A",X"0C",
		X"62",X"D6",X"0E",X"BA",X"D2",X"1B",X"2A",X"3A",X"10",X"62",X"A7",X"3A",X"03",X"62",X"CA",X"08",
		X"2A",X"F6",X"07",X"D6",X"04",X"C3",X"0E",X"2A",X"D6",X"08",X"F6",X"07",X"C6",X"04",X"32",X"03",
		X"62",X"32",X"72",X"69",X"3E",X"01",X"06",X"00",X"33",X"33",X"C9",X"AF",X"32",X"00",X"62",X"C9",
		X"47",X"C9",X"06",X"06",X"11",X"10",X"00",X"DD",X"21",X"00",X"66",X"CD",X"13",X"29",X"C9",X"DD",
		X"7E",X"03",X"67",X"DD",X"7E",X"05",X"C6",X"04",X"6F",X"E5",X"CD",X"F0",X"2F",X"D1",X"7E",X"FE",
		X"B0",X"DA",X"7B",X"2A",X"E6",X"0F",X"FE",X"08",X"D2",X"7B",X"2A",X"7E",X"FE",X"C0",X"CA",X"7B",
		X"2A",X"DA",X"69",X"2A",X"FE",X"D0",X"DA",X"6E",X"2A",X"FE",X"E0",X"DA",X"63",X"2A",X"FE",X"F0",
		X"DA",X"6E",X"2A",X"E6",X"0F",X"3D",X"C3",X"72",X"2A",X"3E",X"FF",X"C3",X"72",X"2A",X"E6",X"0F",
		X"D6",X"09",X"4F",X"7B",X"E6",X"F8",X"81",X"BB",X"DA",X"7D",X"2A",X"AF",X"C9",X"D6",X"04",X"DD",
		X"77",X"05",X"3E",X"01",X"C9",X"3A",X"15",X"62",X"A7",X"C0",X"3A",X"16",X"62",X"A7",X"C0",X"3A",
		X"98",X"63",X"FE",X"01",X"C8",X"3A",X"03",X"62",X"D6",X"03",X"67",X"3A",X"05",X"62",X"C6",X"0C",
		X"6F",X"E5",X"CD",X"F0",X"2F",X"D1",X"7E",X"FE",X"B0",X"DA",X"B4",X"2A",X"E6",X"0F",X"FE",X"08",
		X"D2",X"B4",X"2A",X"C9",X"7A",X"E6",X"07",X"CA",X"CD",X"2A",X"01",X"20",X"00",X"ED",X"42",X"7E",
		X"FE",X"B0",X"DA",X"CD",X"2A",X"E6",X"0F",X"FE",X"08",X"D2",X"CD",X"2A",X"C9",X"3E",X"01",X"32",
		X"21",X"62",X"C9",X"3A",X"03",X"62",X"47",X"3A",X"05",X"62",X"FE",X"50",X"CA",X"EA",X"2A",X"FE",
		X"78",X"CA",X"F6",X"2A",X"FE",X"C8",X"CA",X"F0",X"2A",X"C9",X"3A",X"A3",X"63",X"C3",X"02",X"2B",
		X"3A",X"A6",X"63",X"C3",X"02",X"2B",X"78",X"FE",X"80",X"3A",X"A5",X"63",X"D2",X"02",X"2B",X"3A",
		X"A4",X"63",X"80",X"32",X"03",X"62",X"32",X"72",X"69",X"CD",X"1F",X"24",X"21",X"03",X"62",X"1D",
		X"CA",X"18",X"2B",X"15",X"CA",X"1A",X"2B",X"C9",X"35",X"C9",X"34",X"C9",X"DD",X"21",X"00",X"62",
		X"CD",X"29",X"2B",X"CD",X"AF",X"29",X"AF",X"47",X"C9",X"3A",X"27",X"62",X"3D",X"C2",X"53",X"2B",
		X"3A",X"03",X"62",X"67",X"3A",X"05",X"62",X"C6",X"07",X"6F",X"CD",X"9B",X"2B",X"A7",X"CA",X"51",
		X"2B",X"7B",X"91",X"FE",X"04",X"D2",X"74",X"2B",X"79",X"D6",X"07",X"32",X"05",X"62",X"3E",X"01",
		X"47",X"E1",X"C9",X"3A",X"03",X"62",X"D6",X"03",X"67",X"3A",X"05",X"62",X"C6",X"07",X"6F",X"CD",
		X"9B",X"2B",X"FE",X"02",X"CA",X"7A",X"2B",X"7A",X"C6",X"07",X"67",X"6B",X"CD",X"9B",X"2B",X"A7",
		X"C8",X"C3",X"7A",X"2B",X"3E",X"00",X"06",X"00",X"E1",X"C9",X"3A",X"10",X"62",X"A7",X"3A",X"03",
		X"62",X"CA",X"8B",X"2B",X"F6",X"07",X"D6",X"04",X"C3",X"91",X"2B",X"D6",X"08",X"F6",X"07",X"C6",
		X"04",X"32",X"03",X"62",X"32",X"70",X"69",X"3E",X"01",X"E1",X"C9",X"E5",X"CD",X"F0",X"2F",X"D1",
		X"7E",X"FE",X"B0",X"DA",X"D9",X"2B",X"E6",X"0F",X"FE",X"08",X"D2",X"D9",X"2B",X"7E",X"FE",X"C0",
		X"CA",X"D9",X"2B",X"DA",X"DC",X"2B",X"FE",X"D0",X"DA",X"CB",X"2B",X"FE",X"E0",X"DA",X"C5",X"2B",
		X"FE",X"F0",X"DA",X"CB",X"2B",X"E6",X"0F",X"3D",X"C3",X"CF",X"2B",X"E6",X"0F",X"D6",X"09",X"4F",
		X"7B",X"E6",X"F8",X"81",X"4F",X"BB",X"DA",X"E1",X"2B",X"AF",X"47",X"C9",X"7B",X"E6",X"F8",X"3D",
		X"4F",X"3A",X"0C",X"62",X"DD",X"96",X"05",X"83",X"B9",X"CA",X"EF",X"2B",X"D2",X"F8",X"2B",X"79",
		X"D6",X"07",X"32",X"05",X"62",X"C3",X"FD",X"2B",X"3E",X"02",X"06",X"00",X"C9",X"3E",X"01",X"47",
		X"E1",X"E1",X"C9",X"3E",X"01",X"F7",X"D7",X"3A",X"93",X"63",X"0F",X"D8",X"3A",X"B1",X"62",X"A7",
		X"C8",X"4F",X"3A",X"B0",X"62",X"D6",X"02",X"B9",X"DA",X"7B",X"2C",X"3A",X"82",X"63",X"CB",X"4F",
		X"C2",X"86",X"2C",X"3A",X"80",X"63",X"47",X"3A",X"1A",X"60",X"E6",X"1F",X"B8",X"CA",X"33",X"2C",
		X"10",X"FA",X"C9",X"3A",X"B0",X"62",X"CB",X"3F",X"B9",X"DA",X"41",X"2C",X"3A",X"19",X"60",X"0F",
		X"D0",X"CD",X"57",X"00",X"E6",X"0F",X"C2",X"86",X"2C",X"3E",X"01",X"32",X"82",X"63",X"3C",X"32",
		X"8F",X"63",X"3E",X"01",X"32",X"92",X"63",X"3A",X"B2",X"62",X"B9",X"C0",X"D6",X"08",X"32",X"B2",
		X"62",X"11",X"20",X"00",X"21",X"00",X"64",X"06",X"05",X"7E",X"A7",X"CA",X"72",X"2C",X"19",X"10",
		X"F8",X"C9",X"3A",X"82",X"63",X"F6",X"80",X"32",X"82",X"63",X"C9",X"C6",X"02",X"B9",X"CA",X"49",
		X"2C",X"3E",X"02",X"C3",X"4B",X"2C",X"AF",X"32",X"82",X"63",X"3E",X"03",X"C3",X"4F",X"2C",X"3E",
		X"01",X"F7",X"D7",X"3A",X"93",X"63",X"0F",X"DA",X"15",X"2D",X"3A",X"92",X"63",X"0F",X"D0",X"DD",
		X"21",X"00",X"67",X"11",X"20",X"00",X"06",X"04",X"DD",X"7E",X"00",X"0F",X"DA",X"B3",X"2C",X"0F",
		X"D2",X"B8",X"2C",X"DD",X"19",X"10",X"F1",X"C9",X"DD",X"22",X"AA",X"62",X"DD",X"36",X"00",X"02",
		X"16",X"00",X"C3",X"6F",X"3F",X"87",X"87",X"5F",X"21",X"7C",X"69",X"19",X"22",X"AC",X"62",X"3E",
		X"01",X"32",X"93",X"63",X"11",X"01",X"05",X"CD",X"9F",X"30",X"21",X"B1",X"62",X"35",X"C2",X"E6",
		X"2C",X"3E",X"01",X"32",X"86",X"63",X"7E",X"FE",X"04",X"D2",X"F6",X"2C",X"21",X"A8",X"69",X"87",
		X"87",X"5F",X"16",X"00",X"19",X"72",X"DD",X"36",X"07",X"15",X"DD",X"36",X"08",X"18",X"DD",X"36",
		X"15",X"00",X"3A",X"82",X"63",X"07",X"D2",X"15",X"2D",X"DD",X"36",X"07",X"19",X"DD",X"36",X"08",
		X"18",X"DD",X"36",X"15",X"01",X"21",X"AF",X"62",X"35",X"C0",X"36",X"18",X"3A",X"8F",X"63",X"A7",
		X"CA",X"51",X"2D",X"4F",X"21",X"32",X"39",X"3A",X"82",X"63",X"0F",X"DA",X"2F",X"2D",X"0D",X"79",
		X"87",X"87",X"87",X"4F",X"87",X"87",X"81",X"5F",X"16",X"00",X"19",X"CD",X"4E",X"00",X"21",X"8F",
		X"63",X"35",X"C2",X"51",X"2D",X"3E",X"01",X"32",X"AF",X"62",X"3A",X"82",X"63",X"0F",X"DA",X"83",
		X"2D",X"2A",X"A8",X"62",X"7E",X"DD",X"2A",X"AA",X"62",X"ED",X"5B",X"AC",X"62",X"FE",X"7F",X"CA",
		X"8C",X"2D",X"4F",X"E6",X"7F",X"12",X"DD",X"7E",X"07",X"CB",X"79",X"CA",X"70",X"2D",X"EE",X"03",
		X"13",X"12",X"DD",X"77",X"07",X"DD",X"7E",X"08",X"13",X"12",X"23",X"7E",X"13",X"12",X"23",X"22",
		X"A8",X"62",X"C9",X"21",X"CC",X"39",X"22",X"A8",X"62",X"C3",X"54",X"2D",X"21",X"C3",X"39",X"22",
		X"A8",X"62",X"DD",X"36",X"01",X"01",X"3A",X"82",X"63",X"0F",X"DA",X"A5",X"2D",X"DD",X"36",X"01",
		X"00",X"DD",X"36",X"02",X"02",X"DD",X"36",X"00",X"01",X"DD",X"36",X"0F",X"01",X"AF",X"DD",X"77",
		X"10",X"DD",X"77",X"11",X"DD",X"77",X"12",X"DD",X"77",X"13",X"DD",X"77",X"14",X"32",X"93",X"63",
		X"32",X"92",X"63",X"1A",X"DD",X"77",X"03",X"13",X"13",X"13",X"1A",X"DD",X"77",X"05",X"21",X"5C",
		X"38",X"CD",X"4E",X"00",X"21",X"0B",X"69",X"0E",X"FC",X"FF",X"C9",X"3E",X"0A",X"F7",X"D7",X"3A",
		X"80",X"63",X"3C",X"A7",X"1F",X"47",X"3A",X"27",X"62",X"FE",X"02",X"20",X"01",X"04",X"3E",X"FE",
		X"37",X"1F",X"A7",X"10",X"FC",X"47",X"3A",X"1A",X"60",X"A0",X"C0",X"3E",X"01",X"32",X"A0",X"63",
		X"32",X"9A",X"63",X"C9",X"3E",X"04",X"F7",X"D7",X"DD",X"21",X"00",X"65",X"FD",X"21",X"7C",X"69",
		X"06",X"02",X"DD",X"7E",X"00",X"0F",X"D2",X"A7",X"2E",X"3A",X"1A",X"60",X"E6",X"0F",X"C2",X"29",
		X"2E",X"FD",X"7E",X"00",X"EE",X"07",X"FD",X"77",X"00",X"DD",X"7E",X"0D",X"FE",X"04",X"CA",X"84",
		X"2E",X"DD",X"34",X"03",X"DD",X"34",X"03",X"DD",X"6E",X"0E",X"DD",X"66",X"0F",X"7E",X"4F",X"FE",
		X"7F",X"CA",X"9C",X"2E",X"23",X"DD",X"86",X"05",X"DD",X"77",X"05",X"DD",X"75",X"0E",X"DD",X"74",
		X"0F",X"DD",X"7E",X"03",X"FE",X"B7",X"DA",X"6C",X"2E",X"79",X"FE",X"7F",X"C2",X"6C",X"2E",X"DD",
		X"36",X"0D",X"04",X"AF",X"32",X"83",X"60",X"3E",X"03",X"32",X"84",X"60",X"DD",X"7E",X"03",X"FD",
		X"77",X"02",X"DD",X"7E",X"05",X"FD",X"77",X"03",X"11",X"10",X"00",X"DD",X"19",X"1E",X"04",X"FD",
		X"19",X"10",X"8F",X"C9",X"3E",X"03",X"DD",X"86",X"05",X"DD",X"77",X"05",X"FE",X"F8",X"DA",X"6C",
		X"2E",X"DD",X"36",X"03",X"00",X"DD",X"36",X"00",X"00",X"C3",X"6C",X"2E",X"21",X"AA",X"39",X"3E",
		X"03",X"32",X"83",X"60",X"C3",X"4B",X"2E",X"3A",X"96",X"63",X"0F",X"D2",X"78",X"2E",X"AF",X"32",
		X"96",X"63",X"DD",X"36",X"05",X"50",X"DD",X"36",X"0D",X"01",X"CD",X"57",X"00",X"E6",X"0F",X"C6",
		X"F8",X"DD",X"77",X"03",X"DD",X"36",X"00",X"01",X"21",X"AA",X"39",X"DD",X"75",X"0E",X"DD",X"74",
		X"0F",X"C3",X"78",X"2E",X"3E",X"0B",X"F7",X"D7",X"11",X"8C",X"69",X"DD",X"21",X"80",X"66",X"DD",
		X"7E",X"01",X"0F",X"DA",X"ED",X"2E",X"00",X"00",X"00",X"DD",X"21",X"90",X"66",X"DD",X"36",X"0E",
		X"00",X"DD",X"36",X"0F",X"F0",X"3A",X"17",X"62",X"0F",X"D2",X"97",X"2F",X"AF",X"32",X"18",X"62",
		X"21",X"89",X"60",X"00",X"00",X"DD",X"36",X"09",X"06",X"DD",X"36",X"0A",X"03",X"06",X"1E",X"3A",
		X"07",X"62",X"CB",X"27",X"D2",X"1B",X"2F",X"F6",X"80",X"CB",X"F8",X"F6",X"08",X"4F",X"3A",X"94",
		X"63",X"CB",X"5F",X"CA",X"43",X"2F",X"CB",X"C0",X"CB",X"C1",X"DD",X"36",X"09",X"05",X"DD",X"36",
		X"0A",X"06",X"DD",X"36",X"0F",X"00",X"DD",X"36",X"0E",X"F0",X"CB",X"79",X"CA",X"43",X"2F",X"DD",
		X"36",X"0E",X"10",X"79",X"32",X"70",X"69",X"0E",X"10",X"21",X"94",X"63",X"34",X"C2",X"B7",X"2F",
		X"21",X"95",X"63",X"34",X"7E",X"FE",X"02",X"C2",X"BE",X"2F",X"AF",X"32",X"95",X"63",X"32",X"17",
		X"62",X"DD",X"77",X"01",X"3A",X"03",X"62",X"ED",X"44",X"DD",X"77",X"0E",X"3A",X"07",X"62",X"32",
		X"70",X"69",X"DD",X"36",X"00",X"00",X"3A",X"89",X"63",X"32",X"89",X"60",X"EB",X"3A",X"03",X"62",
		X"DD",X"86",X"0E",X"DD",X"77",X"03",X"2C",X"2C",X"77",X"2B",X"2B",X"70",X"2C",X"71",X"2C",X"2C",
		X"3A",X"05",X"62",X"C3",X"3B",X"3F",X"C9",X"3A",X"18",X"62",X"0F",X"D0",X"DD",X"36",X"09",X"06",
		X"DD",X"36",X"0A",X"03",X"3A",X"07",X"62",X"07",X"3E",X"3C",X"1F",X"47",X"0E",X"10",X"3A",X"89",
		X"60",X"32",X"89",X"63",X"C3",X"7C",X"2F",X"3A",X"95",X"63",X"A7",X"CA",X"7C",X"2F",X"3A",X"1A",
		X"60",X"CB",X"5F",X"CA",X"7C",X"2F",X"0E",X"10",X"C3",X"7C",X"2F",X"3E",X"0E",X"F7",X"21",X"B4",
		X"62",X"35",X"C0",X"3E",X"03",X"32",X"B9",X"62",X"32",X"96",X"63",X"11",X"01",X"05",X"CD",X"9F",
		X"30",X"3A",X"B3",X"62",X"77",X"21",X"B1",X"62",X"35",X"C0",X"3E",X"01",X"32",X"86",X"63",X"C9",
		X"7D",X"0F",X"0F",X"0F",X"E6",X"1F",X"6F",X"7C",X"2F",X"E6",X"F8",X"5F",X"AF",X"67",X"CB",X"13",
		X"17",X"CB",X"13",X"17",X"C6",X"90",X"57",X"19",X"C9",X"57",X"0F",X"DA",X"22",X"30",X"0E",X"93",
		X"0F",X"0F",X"D2",X"17",X"30",X"0E",X"6C",X"07",X"DA",X"31",X"30",X"79",X"E6",X"F0",X"4F",X"C3",
		X"31",X"30",X"0E",X"B4",X"0F",X"0F",X"D2",X"2B",X"30",X"0E",X"1E",X"CB",X"50",X"CA",X"31",X"30",
		X"05",X"79",X"0F",X"0F",X"4F",X"E6",X"03",X"B8",X"C2",X"31",X"30",X"79",X"0F",X"0F",X"E6",X"03",
		X"FE",X"03",X"C0",X"CB",X"92",X"15",X"C0",X"3E",X"04",X"C9",X"11",X"E0",X"FF",X"3A",X"8E",X"63",
		X"4F",X"06",X"00",X"21",X"00",X"92",X"CD",X"64",X"30",X"21",X"C0",X"91",X"CD",X"64",X"30",X"21",
		X"8E",X"63",X"35",X"C9",X"09",X"7E",X"19",X"77",X"C9",X"DF",X"2A",X"C0",X"63",X"34",X"C9",X"21",
		X"AF",X"62",X"34",X"7E",X"E6",X"07",X"C0",X"21",X"73",X"69",X"0E",X"FC",X"FF",X"0E",X"81",X"21",
		X"70",X"69",X"CD",X"96",X"30",X"21",X"84",X"69",X"CD",X"96",X"30",X"CD",X"57",X"00",X"E6",X"80",
		X"00",X"00",X"00",X"AE",X"77",X"C9",X"06",X"02",X"79",X"AE",X"77",X"19",X"10",X"FA",X"C9",X"E5",
		X"21",X"C0",X"60",X"3A",X"B0",X"60",X"6F",X"CB",X"7E",X"CA",X"BB",X"30",X"72",X"2C",X"73",X"2C",
		X"7D",X"FE",X"C0",X"D2",X"B8",X"30",X"3E",X"C0",X"32",X"B0",X"60",X"E1",X"C9",X"21",X"50",X"69",
		X"06",X"02",X"00",X"00",X"00",X"2E",X"80",X"06",X"0A",X"00",X"00",X"00",X"2E",X"B8",X"06",X"0B",
		X"00",X"00",X"00",X"21",X"0C",X"6A",X"06",X"05",X"C3",X"E4",X"30",X"CD",X"11",X"4C",X"C9",X"00",
		X"2E",X"58",X"06",X"06",X"7D",X"36",X"3F",X"C6",X"04",X"6F",X"10",X"F9",X"C9",X"CD",X"FA",X"30",
		X"CD",X"3C",X"31",X"CD",X"B1",X"31",X"CD",X"F3",X"34",X"C9",X"3A",X"80",X"63",X"FE",X"06",X"38",
		X"02",X"3E",X"05",X"EF",X"10",X"31",X"10",X"31",X"1B",X"31",X"26",X"31",X"26",X"31",X"31",X"31",
		X"3A",X"1A",X"60",X"E6",X"01",X"FE",X"01",X"C8",X"33",X"33",X"C9",X"3A",X"1A",X"60",X"E6",X"07",
		X"FE",X"05",X"F8",X"33",X"33",X"C9",X"3A",X"1A",X"60",X"E6",X"03",X"FE",X"03",X"F8",X"33",X"33",
		X"C9",X"3A",X"1A",X"60",X"E6",X"07",X"FE",X"07",X"F8",X"33",X"33",X"C9",X"DD",X"21",X"00",X"64",
		X"AF",X"32",X"A1",X"63",X"00",X"00",X"CD",X"E3",X"42",X"DD",X"7E",X"00",X"FE",X"00",X"CA",X"7C",
		X"31",X"3A",X"A1",X"63",X"3C",X"32",X"A1",X"63",X"3E",X"1E",X"DD",X"77",X"08",X"3A",X"17",X"62",
		X"FE",X"01",X"C2",X"6A",X"31",X"3E",X"1D",X"DD",X"77",X"08",X"DD",X"19",X"10",X"DB",X"21",X"A0",
		X"63",X"36",X"00",X"3A",X"A1",X"63",X"FE",X"00",X"C0",X"33",X"33",X"C9",X"3A",X"A1",X"63",X"FE",
		X"05",X"CA",X"6A",X"31",X"3A",X"27",X"62",X"FE",X"02",X"C2",X"95",X"31",X"3A",X"A1",X"63",X"4F",
		X"3A",X"80",X"63",X"B9",X"C8",X"3A",X"A0",X"63",X"FE",X"01",X"C2",X"6A",X"31",X"DD",X"77",X"00",
		X"DD",X"77",X"18",X"AF",X"32",X"A0",X"63",X"3A",X"A1",X"63",X"3C",X"32",X"A1",X"63",X"C3",X"6A",
		X"31",X"CD",X"DD",X"31",X"AF",X"32",X"A2",X"63",X"21",X"E0",X"63",X"22",X"C8",X"63",X"2A",X"C8",
		X"63",X"01",X"20",X"00",X"09",X"22",X"C8",X"63",X"7E",X"A7",X"CA",X"D0",X"31",X"CD",X"02",X"32",
		X"3A",X"A2",X"63",X"3C",X"32",X"A2",X"63",X"FE",X"05",X"C2",X"BE",X"31",X"C9",X"3A",X"80",X"63",
		X"FE",X"03",X"F8",X"CD",X"F6",X"31",X"FE",X"01",X"C0",X"21",X"39",X"64",X"3E",X"02",X"77",X"21",
		X"79",X"64",X"3E",X"02",X"77",X"C9",X"3A",X"18",X"60",X"E6",X"03",X"FE",X"01",X"C0",X"3A",X"1A",
		X"60",X"C9",X"DD",X"2A",X"C8",X"63",X"DD",X"7E",X"18",X"FE",X"01",X"CA",X"7A",X"32",X"DD",X"7E",
		X"0D",X"FE",X"04",X"F2",X"30",X"32",X"DD",X"7E",X"19",X"FE",X"02",X"CA",X"7E",X"32",X"CD",X"0F",
		X"33",X"3A",X"18",X"60",X"E6",X"03",X"C2",X"33",X"32",X"DD",X"7E",X"0D",X"A7",X"CA",X"57",X"32",
		X"CD",X"3D",X"33",X"DD",X"7E",X"0D",X"FE",X"04",X"F2",X"91",X"32",X"CD",X"AD",X"33",X"CD",X"8C",
		X"29",X"FE",X"01",X"CA",X"97",X"32",X"DD",X"2A",X"C8",X"63",X"DD",X"7E",X"0E",X"FE",X"10",X"DA",
		X"8C",X"32",X"FE",X"F0",X"D2",X"84",X"32",X"DD",X"7E",X"13",X"FE",X"00",X"C2",X"B9",X"32",X"3E",
		X"11",X"DD",X"77",X"13",X"16",X"00",X"5F",X"21",X"7A",X"3A",X"19",X"7E",X"DD",X"46",X"0E",X"DD",
		X"70",X"03",X"DD",X"4E",X"0F",X"81",X"DD",X"77",X"05",X"C9",X"CD",X"BD",X"32",X"C9",X"CD",X"D6",
		X"32",X"C3",X"29",X"32",X"3E",X"02",X"DD",X"77",X"0D",X"C3",X"57",X"32",X"3E",X"01",X"C3",X"86",
		X"32",X"CD",X"E7",X"33",X"C3",X"57",X"32",X"DD",X"2A",X"C8",X"63",X"DD",X"7E",X"0D",X"FE",X"01",
		X"C2",X"B1",X"32",X"3E",X"02",X"DD",X"35",X"0E",X"DD",X"77",X"0D",X"CD",X"C3",X"33",X"C3",X"57",
		X"32",X"3E",X"01",X"DD",X"34",X"0E",X"C3",X"A8",X"32",X"3D",X"C3",X"61",X"32",X"3A",X"27",X"62",
		X"FE",X"01",X"CA",X"CE",X"32",X"FE",X"02",X"CA",X"D2",X"32",X"CD",X"B9",X"34",X"C9",X"CD",X"2C",
		X"34",X"C9",X"CD",X"78",X"34",X"C9",X"DD",X"7E",X"1C",X"FE",X"00",X"C2",X"FD",X"32",X"DD",X"7E",
		X"1D",X"FE",X"01",X"C2",X"0B",X"33",X"DD",X"36",X"1D",X"00",X"3A",X"05",X"62",X"DD",X"46",X"0F",
		X"90",X"DA",X"03",X"33",X"DD",X"36",X"1C",X"FF",X"DD",X"36",X"0D",X"00",X"C9",X"DD",X"35",X"1C",
		X"C2",X"F8",X"32",X"DD",X"36",X"19",X"00",X"DD",X"36",X"1C",X"00",X"CD",X"0F",X"33",X"C9",X"DD",
		X"7E",X"16",X"FE",X"00",X"C2",X"32",X"33",X"DD",X"36",X"16",X"2B",X"DD",X"36",X"0D",X"00",X"3A",
		X"18",X"60",X"0F",X"D2",X"32",X"33",X"DD",X"7E",X"0D",X"FE",X"01",X"CA",X"36",X"33",X"DD",X"36",
		X"0D",X"01",X"DD",X"35",X"16",X"C9",X"DD",X"36",X"0D",X"02",X"C3",X"32",X"33",X"DD",X"7E",X"0D",
		X"FE",X"08",X"CA",X"71",X"33",X"FE",X"04",X"CA",X"8A",X"33",X"CD",X"A1",X"33",X"DD",X"7E",X"0F",
		X"C6",X"08",X"57",X"DD",X"7E",X"0E",X"01",X"15",X"00",X"CD",X"6E",X"23",X"A7",X"CA",X"99",X"33",
		X"DD",X"70",X"1F",X"3A",X"05",X"62",X"47",X"DD",X"7E",X"0F",X"90",X"D0",X"DD",X"36",X"0D",X"04",
		X"C9",X"DD",X"7E",X"0F",X"C6",X"08",X"DD",X"46",X"1F",X"B8",X"C0",X"DD",X"36",X"0D",X"00",X"DD",
		X"7E",X"19",X"FE",X"02",X"C0",X"DD",X"36",X"1D",X"01",X"C9",X"DD",X"7E",X"0F",X"C6",X"08",X"DD",
		X"46",X"1F",X"B8",X"C0",X"DD",X"36",X"0D",X"00",X"C9",X"DD",X"70",X"1F",X"DD",X"36",X"0D",X"08",
		X"C9",X"3E",X"07",X"F7",X"DD",X"7E",X"0F",X"FE",X"59",X"D0",X"33",X"33",X"C9",X"DD",X"7E",X"0D",
		X"FE",X"01",X"CA",X"D9",X"33",X"DD",X"7E",X"07",X"E6",X"7F",X"DD",X"77",X"07",X"DD",X"35",X"0E",
		X"CD",X"09",X"34",X"3A",X"27",X"62",X"FE",X"01",X"C0",X"DD",X"66",X"0E",X"DD",X"6E",X"0F",X"DD",
		X"46",X"0D",X"CD",X"33",X"23",X"DD",X"75",X"0F",X"C9",X"DD",X"7E",X"07",X"F6",X"80",X"DD",X"77",
		X"07",X"DD",X"34",X"0E",X"C3",X"C0",X"33",X"CD",X"09",X"34",X"DD",X"7E",X"0D",X"FE",X"08",X"C2",
		X"05",X"34",X"DD",X"7E",X"14",X"A7",X"C2",X"01",X"34",X"DD",X"36",X"14",X"02",X"DD",X"35",X"0F",
		X"C9",X"DD",X"35",X"14",X"C9",X"DD",X"34",X"0F",X"C9",X"DD",X"7E",X"15",X"A7",X"C2",X"28",X"34",
		X"DD",X"36",X"15",X"02",X"DD",X"34",X"07",X"DD",X"7E",X"07",X"E6",X"0F",X"FE",X"0F",X"C0",X"DD",
		X"7E",X"07",X"EE",X"02",X"DD",X"77",X"07",X"C9",X"DD",X"35",X"15",X"C9",X"DD",X"6E",X"1A",X"DD",
		X"66",X"1B",X"AF",X"01",X"00",X"00",X"ED",X"4A",X"C2",X"42",X"34",X"21",X"8C",X"3A",X"DD",X"36",
		X"03",X"26",X"DD",X"34",X"03",X"7E",X"FE",X"AA",X"CA",X"56",X"34",X"DD",X"77",X"05",X"23",X"DD",
		X"75",X"1A",X"DD",X"74",X"1B",X"C9",X"AF",X"DD",X"77",X"13",X"DD",X"77",X"18",X"DD",X"77",X"0D",
		X"DD",X"77",X"1C",X"DD",X"7E",X"03",X"DD",X"77",X"0E",X"DD",X"7E",X"05",X"DD",X"77",X"0F",X"DD",
		X"36",X"1A",X"00",X"DD",X"36",X"1B",X"00",X"C9",X"DD",X"6E",X"1A",X"DD",X"66",X"1B",X"AF",X"01",
		X"00",X"00",X"ED",X"4A",X"C2",X"9A",X"34",X"21",X"AC",X"3A",X"3A",X"03",X"62",X"CB",X"7F",X"CA",
		X"A8",X"34",X"DD",X"36",X"0D",X"01",X"DD",X"36",X"03",X"7E",X"DD",X"7E",X"0D",X"FE",X"01",X"C2",
		X"B3",X"34",X"DD",X"34",X"03",X"C3",X"45",X"34",X"DD",X"36",X"0D",X"02",X"DD",X"36",X"03",X"80",
		X"C3",X"9A",X"34",X"DD",X"35",X"03",X"C3",X"45",X"34",X"3A",X"27",X"62",X"FE",X"03",X"C8",X"3A",
		X"03",X"62",X"CB",X"7F",X"C2",X"ED",X"34",X"21",X"C4",X"3A",X"06",X"00",X"3A",X"19",X"60",X"E6",
		X"06",X"4F",X"09",X"7E",X"DD",X"77",X"03",X"DD",X"77",X"0E",X"23",X"7E",X"DD",X"77",X"05",X"DD",
		X"77",X"0F",X"AF",X"DD",X"77",X"0D",X"DD",X"77",X"18",X"DD",X"77",X"1C",X"C9",X"21",X"D4",X"3A",
		X"C3",X"CA",X"34",X"21",X"00",X"64",X"CD",X"C3",X"42",X"00",X"00",X"7E",X"A7",X"CA",X"1E",X"35",
		X"CD",X"F5",X"42",X"7E",X"12",X"23",X"1C",X"7E",X"12",X"7D",X"D6",X"05",X"6F",X"1C",X"7E",X"12",
		X"00",X"23",X"23",X"1C",X"7E",X"12",X"13",X"3E",X"1B",X"85",X"6F",X"10",X"DE",X"C9",X"3E",X"05",
		X"85",X"6F",X"3E",X"04",X"83",X"5F",X"C3",X"17",X"35",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"02",X"00",X"00",X"03",X"00",X"00",X"04",X"00",X"00",X"05",X"00",X"00",X"06",X"00",X"00",X"07",
		X"00",X"00",X"08",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"20",X"00",
		X"00",X"30",X"00",X"00",X"40",X"00",X"00",X"50",X"00",X"00",X"60",X"00",X"00",X"70",X"00",X"00",
		X"80",X"00",X"00",X"90",X"00",X"94",X"93",X"01",X"23",X"24",X"FD",X"FD",X"00",X"00",X"07",X"06",
		X"05",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"3F",X"00",X"50",X"76",X"00",X"F4",X"76",X"96",X"93",X"02",X"1E",X"14",X"FD",X"FD",X"00",X"00",
		X"06",X"01",X"00",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"3F",X"00",X"00",X"61",X"00",X"F6",X"76",X"98",X"93",X"03",X"22",X"14",X"FD",X"FD",
		X"00",X"00",X"05",X"09",X"05",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"3F",X"00",X"50",X"59",X"00",X"F8",X"76",X"9A",X"93",X"04",X"24",X"18",
		X"FD",X"FD",X"00",X"00",X"05",X"00",X"05",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"3F",X"00",X"50",X"50",X"00",X"FA",X"76",X"9C",X"93",X"05",
		X"24",X"18",X"FD",X"FD",X"00",X"00",X"04",X"03",X"00",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"3F",X"00",X"00",X"43",X"00",X"FC",X"92",X"3B",
		X"5C",X"4B",X"5C",X"5B",X"5C",X"6B",X"5C",X"7B",X"5C",X"8B",X"5C",X"9B",X"5C",X"AB",X"5C",X"BB",
		X"5C",X"CB",X"5C",X"3B",X"6C",X"4B",X"6C",X"5B",X"6C",X"6B",X"6C",X"7B",X"6C",X"8B",X"6C",X"9B",
		X"6C",X"AB",X"6C",X"BB",X"6C",X"CB",X"6C",X"3B",X"7C",X"4B",X"7C",X"5B",X"7C",X"6B",X"7C",X"7B",
		X"7C",X"8B",X"7C",X"9B",X"7C",X"AB",X"7C",X"BB",X"7C",X"CB",X"7C",X"8B",X"36",X"01",X"00",X"98",
		X"36",X"A5",X"36",X"B2",X"36",X"BF",X"36",X"06",X"00",X"CC",X"36",X"08",X"00",X"E6",X"36",X"FD",
		X"36",X"0B",X"00",X"15",X"37",X"1C",X"37",X"30",X"37",X"38",X"37",X"47",X"37",X"5D",X"37",X"73",
		X"37",X"8B",X"37",X"00",X"61",X"22",X"61",X"44",X"61",X"66",X"61",X"88",X"61",X"9E",X"37",X"B6",
		X"37",X"D2",X"37",X"E1",X"37",X"1D",X"00",X"F4",X"37",X"06",X"38",X"96",X"92",X"17",X"11",X"1D",
		X"15",X"FD",X"FD",X"1F",X"26",X"15",X"22",X"3F",X"94",X"92",X"20",X"1C",X"11",X"29",X"15",X"22",
		X"FD",X"30",X"32",X"31",X"3F",X"94",X"92",X"20",X"1C",X"11",X"29",X"15",X"22",X"FD",X"30",X"33",
		X"31",X"3F",X"80",X"92",X"18",X"19",X"17",X"18",X"FD",X"23",X"13",X"1F",X"22",X"15",X"3F",X"9F",
		X"91",X"13",X"22",X"15",X"14",X"19",X"24",X"FD",X"FD",X"FD",X"FD",X"3F",X"5E",X"93",X"18",X"1F",
		X"27",X"FD",X"18",X"19",X"17",X"18",X"FD",X"13",X"11",X"1E",X"FD",X"29",X"1F",X"25",X"FD",X"24",
		X"22",X"29",X"FD",X"FB",X"FD",X"3F",X"29",X"93",X"1F",X"1E",X"1C",X"29",X"FD",X"01",X"FD",X"20",
		X"1C",X"11",X"29",X"15",X"22",X"FD",X"12",X"25",X"24",X"24",X"1F",X"1E",X"3F",X"29",X"93",X"01",
		X"FD",X"1F",X"22",X"FD",X"02",X"FD",X"20",X"1C",X"11",X"29",X"15",X"22",X"23",X"FD",X"12",X"25",
		X"24",X"24",X"1F",X"1E",X"3F",X"27",X"92",X"20",X"25",X"23",X"18",X"3F",X"06",X"93",X"1E",X"11",
		X"1D",X"15",X"FD",X"22",X"15",X"17",X"19",X"23",X"24",X"22",X"11",X"24",X"19",X"1F",X"1E",X"3F",
		X"88",X"92",X"1E",X"11",X"1D",X"15",X"2E",X"3F",X"E9",X"75",X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"3F",X"0B",X"93",X"11",X"FD",X"12",X"FD",X"13",X"FD",X"14",
		X"FD",X"15",X"FD",X"16",X"FD",X"17",X"FD",X"18",X"FD",X"19",X"FD",X"1A",X"3F",X"0D",X"93",X"1B",
		X"FD",X"1C",X"FD",X"1D",X"FD",X"1E",X"FD",X"1F",X"FD",X"20",X"FD",X"21",X"FD",X"22",X"FD",X"23",
		X"FD",X"24",X"3F",X"0F",X"93",X"25",X"FD",X"26",X"FD",X"27",X"FD",X"28",X"FD",X"29",X"FD",X"2A",
		X"FD",X"2B",X"FD",X"2C",X"44",X"45",X"46",X"47",X"48",X"FD",X"3F",X"F2",X"92",X"22",X"15",X"17",
		X"19",X"FD",X"24",X"19",X"1D",X"15",X"FD",X"FD",X"30",X"06",X"00",X"31",X"FD",X"3F",X"92",X"93",
		X"22",X"11",X"1E",X"1B",X"FD",X"FD",X"23",X"13",X"1F",X"22",X"15",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"FD",X"1E",X"11",X"1D",X"15",X"3F",X"72",X"93",X"29",X"1F",X"25",X"22",X"FD",X"1E",X"11",X"1D",
		X"15",X"FD",X"27",X"11",X"23",X"FD",X"22",X"15",X"17",X"19",X"23",X"24",X"15",X"22",X"15",X"14",
		X"42",X"3F",X"A7",X"92",X"19",X"1E",X"23",X"15",X"22",X"24",X"FD",X"13",X"1F",X"19",X"1E",X"FD",
		X"3F",X"0A",X"93",X"FD",X"FD",X"20",X"1C",X"11",X"29",X"15",X"22",X"FD",X"FD",X"FD",X"FD",X"13",
		X"1F",X"19",X"1E",X"3F",X"0C",X"90",X"49",X"4A",X"FD",X"1E",X"19",X"1E",X"24",X"15",X"1E",X"14",
		X"1F",X"FD",X"FD",X"FD",X"FD",X"3F",X"BD",X"91",X"01",X"09",X"08",X"01",X"3F",X"02",X"97",X"38",
		X"68",X"38",X"02",X"DF",X"54",X"10",X"54",X"02",X"EF",X"6D",X"20",X"6D",X"02",X"DF",X"8E",X"10",
		X"8E",X"02",X"EF",X"AF",X"20",X"AF",X"02",X"DF",X"D0",X"10",X"D0",X"02",X"EF",X"F1",X"10",X"F1",
		X"00",X"53",X"18",X"53",X"54",X"00",X"63",X"18",X"63",X"54",X"00",X"93",X"38",X"93",X"54",X"00",
		X"83",X"54",X"83",X"F1",X"00",X"93",X"54",X"93",X"F1",X"AA",X"8D",X"7D",X"8C",X"6F",X"00",X"7C",
		X"6E",X"00",X"7C",X"6D",X"00",X"7C",X"6C",X"00",X"7C",X"8F",X"7F",X"8E",X"27",X"13",X"47",X"50",
		X"A7",X"13",X"2F",X"50",X"25",X"13",X"3B",X"50",X"3F",X"13",X"00",X"00",X"23",X"13",X"3B",X"40",
		X"A9",X"13",X"46",X"44",X"3F",X"13",X"00",X"00",X"29",X"13",X"30",X"44",X"3F",X"13",X"00",X"48",
		X"70",X"13",X"00",X"48",X"10",X"13",X"6F",X"23",X"11",X"13",X"6F",X"33",X"34",X"13",X"51",X"3C",
		X"35",X"13",X"00",X"3C",X"32",X"13",X"54",X"40",X"33",X"13",X"63",X"40",X"14",X"11",X"6A",X"48",
		X"36",X"13",X"53",X"50",X"37",X"13",X"63",X"50",X"31",X"13",X"6B",X"41",X"3F",X"13",X"6A",X"48",
		X"14",X"11",X"6A",X"48",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"FE",X"FE",X"FE",X"FE",X"FE",
		X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"01",X"01",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"7F",X"04",X"7F",X"F0",X"10",
		X"F0",X"02",X"DF",X"F2",X"70",X"F8",X"02",X"6F",X"F8",X"10",X"F8",X"AA",X"04",X"DF",X"D0",X"90",
		X"D0",X"02",X"DF",X"DC",X"20",X"D1",X"AA",X"FF",X"FF",X"FF",X"FF",X"FF",X"04",X"DF",X"A8",X"20",
		X"A8",X"04",X"5F",X"B0",X"20",X"B0",X"02",X"DF",X"B0",X"20",X"BB",X"AA",X"04",X"DF",X"88",X"30",
		X"88",X"04",X"DF",X"90",X"B0",X"90",X"02",X"DF",X"9A",X"20",X"8F",X"AA",X"04",X"BF",X"68",X"20",
		X"68",X"04",X"3F",X"70",X"20",X"70",X"02",X"DF",X"6E",X"20",X"79",X"AA",X"02",X"DF",X"58",X"A0",
		X"55",X"AA",X"70",X"13",X"00",X"44",X"AC",X"13",X"2B",X"4C",X"AE",X"13",X"3B",X"4C",X"AF",X"13",
		X"3B",X"3C",X"B0",X"13",X"4B",X"3C",X"AD",X"13",X"4B",X"4C",X"70",X"13",X"00",X"44",X"70",X"13",
		X"00",X"44",X"70",X"13",X"00",X"44",X"70",X"13",X"00",X"44",X"27",X"13",X"47",X"4C",X"A7",X"13",
		X"2F",X"4C",X"25",X"13",X"3B",X"4C",X"70",X"13",X"00",X"44",X"23",X"13",X"3B",X"3C",X"2A",X"13",
		X"4B",X"3C",X"2B",X"13",X"4B",X"4C",X"AA",X"18",X"2B",X"3C",X"AB",X"18",X"2B",X"4C",X"70",X"1A",
		X"00",X"44",X"70",X"18",X"00",X"44",X"08",X"18",X"4B",X"4C",X"2E",X"18",X"3B",X"4C",X"08",X"18",
		X"3A",X"3C",X"30",X"17",X"2B",X"3C",X"2D",X"18",X"2B",X"4C",X"70",X"18",X"00",X"44",X"70",X"18",
		X"00",X"44",X"70",X"18",X"00",X"44",X"70",X"1A",X"00",X"44",X"FD",X"FD",X"FD",X"FE",X"FE",X"FE",
		X"FE",X"FF",X"FF",X"00",X"FF",X"00",X"00",X"01",X"00",X"01",X"01",X"02",X"02",X"02",X"02",X"03",
		X"03",X"03",X"7F",X"1E",X"4E",X"BB",X"4C",X"D8",X"4E",X"59",X"4E",X"7F",X"BB",X"4D",X"7F",X"27",
		X"13",X"47",X"50",X"26",X"13",X"2D",X"50",X"25",X"13",X"3B",X"50",X"3F",X"13",X"00",X"48",X"24",
		X"13",X"3B",X"40",X"28",X"13",X"4B",X"40",X"3F",X"13",X"00",X"48",X"29",X"13",X"30",X"44",X"3F",
		X"13",X"00",X"48",X"3F",X"13",X"00",X"48",X"A6",X"13",X"49",X"50",X"A7",X"13",X"2F",X"50",X"25",
		X"13",X"3B",X"50",X"3F",X"13",X"08",X"48",X"24",X"13",X"3B",X"40",X"A9",X"13",X"46",X"44",X"3F",
		X"13",X"00",X"48",X"A8",X"13",X"2B",X"40",X"3F",X"13",X"00",X"48",X"3F",X"13",X"00",X"48",X"E7",
		X"13",X"73",X"60",X"67",X"13",X"8B",X"60",X"65",X"13",X"7F",X"60",X"3F",X"13",X"00",X"68",X"64",
		X"13",X"7F",X"70",X"69",X"13",X"74",X"6C",X"3F",X"13",X"00",X"68",X"E9",X"13",X"8A",X"6C",X"3F",
		X"13",X"00",X"68",X"3F",X"13",X"00",X"68",X"05",X"AF",X"F0",X"50",X"F0",X"AA",X"05",X"AF",X"E8",
		X"50",X"E8",X"AA",X"05",X"AF",X"E0",X"50",X"E0",X"AA",X"05",X"AF",X"D8",X"50",X"D8",X"AA",X"05",
		X"B7",X"58",X"48",X"58",X"AA",X"01",X"02",X"03",X"04",X"01",X"02",X"03",X"04",X"01",X"02",X"03",
		X"04",X"01",X"02",X"03",X"04",X"01",X"02",X"03",X"04",X"7F",X"FF",X"00",X"FF",X"FF",X"FE",X"FE",
		X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"00",X"E8",X"E5",X"E3",X"E2",
		X"E1",X"E0",X"DF",X"DE",X"DD",X"DD",X"DC",X"DC",X"DC",X"DC",X"DC",X"DC",X"DD",X"DD",X"DE",X"DF",
		X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E7",X"E9",X"EB",X"ED",X"F0",X"AA",X"80",X"7B",X"78",X"76",
		X"74",X"73",X"72",X"71",X"70",X"70",X"6F",X"6F",X"6F",X"70",X"70",X"71",X"72",X"73",X"74",X"75",
		X"76",X"77",X"78",X"AA",X"EE",X"F0",X"DB",X"A0",X"E6",X"C8",X"D6",X"78",X"EB",X"F0",X"DB",X"A0",
		X"E6",X"C8",X"E6",X"C8",X"1B",X"C8",X"23",X"A0",X"2B",X"78",X"12",X"F0",X"1B",X"C8",X"23",X"A0",
		X"12",X"F0",X"1B",X"C8",X"02",X"97",X"38",X"68",X"38",X"02",X"9F",X"54",X"10",X"54",X"02",X"DF",
		X"58",X"A0",X"55",X"02",X"EF",X"6D",X"20",X"79",X"02",X"DF",X"9A",X"10",X"8E",X"02",X"EF",X"AF",
		X"20",X"BB",X"02",X"DF",X"DC",X"10",X"D0",X"02",X"FF",X"F0",X"80",X"F7",X"02",X"7F",X"F8",X"00",
		X"F8",X"00",X"CB",X"57",X"CB",X"6F",X"00",X"CB",X"99",X"CB",X"B1",X"00",X"CB",X"DB",X"CB",X"F3",
		X"00",X"63",X"18",X"63",X"54",X"01",X"63",X"D5",X"63",X"F8",X"00",X"33",X"78",X"33",X"90",X"00",
		X"33",X"BA",X"33",X"D2",X"00",X"53",X"18",X"53",X"54",X"01",X"53",X"92",X"53",X"B8",X"00",X"5B",
		X"76",X"5B",X"92",X"00",X"73",X"B6",X"73",X"D6",X"00",X"83",X"95",X"83",X"B5",X"00",X"93",X"38",
		X"93",X"54",X"01",X"BB",X"70",X"BB",X"98",X"01",X"6B",X"54",X"6B",X"75",X"AA",X"06",X"8F",X"90",
		X"70",X"90",X"06",X"8F",X"98",X"70",X"98",X"06",X"8F",X"A0",X"70",X"A0",X"00",X"63",X"18",X"63",
		X"58",X"00",X"63",X"80",X"63",X"A8",X"00",X"63",X"D0",X"63",X"F8",X"00",X"53",X"18",X"53",X"58",
		X"00",X"53",X"A8",X"53",X"D0",X"00",X"9B",X"80",X"9B",X"A8",X"00",X"9B",X"D0",X"9B",X"F8",X"01",
		X"23",X"58",X"23",X"80",X"01",X"DB",X"58",X"DB",X"80",X"00",X"2B",X"80",X"2B",X"A8",X"00",X"D3",
		X"80",X"D3",X"A8",X"00",X"A3",X"A8",X"A3",X"D0",X"00",X"2B",X"D0",X"2B",X"F8",X"00",X"D3",X"D0",
		X"D3",X"F8",X"00",X"93",X"38",X"93",X"58",X"02",X"97",X"38",X"68",X"38",X"03",X"EF",X"58",X"10",
		X"58",X"03",X"F7",X"80",X"88",X"80",X"03",X"77",X"80",X"08",X"80",X"02",X"A7",X"A8",X"50",X"A8",
		X"02",X"E7",X"A8",X"B8",X"A8",X"02",X"3F",X"A8",X"18",X"A8",X"03",X"EF",X"D0",X"10",X"D0",X"02",
		X"EF",X"F8",X"10",X"F8",X"AA",X"00",X"63",X"18",X"63",X"58",X"00",X"63",X"88",X"63",X"D0",X"00",
		X"53",X"18",X"53",X"58",X"00",X"53",X"88",X"53",X"D0",X"00",X"E3",X"68",X"E3",X"90",X"00",X"E3",
		X"B8",X"E3",X"D0",X"00",X"CB",X"90",X"CB",X"B0",X"00",X"B3",X"58",X"B3",X"78",X"00",X"9B",X"80",
		X"9B",X"A0",X"00",X"93",X"38",X"93",X"58",X"00",X"23",X"88",X"23",X"C0",X"00",X"1B",X"C0",X"1B",
		X"E8",X"02",X"97",X"38",X"68",X"38",X"02",X"B7",X"58",X"10",X"58",X"02",X"EF",X"68",X"E0",X"68",
		X"02",X"D7",X"70",X"C8",X"70",X"02",X"BF",X"78",X"B0",X"78",X"02",X"A7",X"80",X"90",X"80",X"02",
		X"67",X"88",X"48",X"88",X"02",X"27",X"88",X"10",X"88",X"02",X"EF",X"90",X"C8",X"90",X"02",X"A7",
		X"A0",X"98",X"A0",X"02",X"BF",X"A8",X"B0",X"A8",X"02",X"D7",X"B0",X"C8",X"B0",X"02",X"EF",X"B8",
		X"E0",X"B8",X"02",X"27",X"C0",X"10",X"C0",X"02",X"EF",X"D0",X"D8",X"D0",X"02",X"67",X"D0",X"50",
		X"D0",X"02",X"CF",X"D8",X"C0",X"D8",X"02",X"B7",X"E0",X"A8",X"E0",X"02",X"9F",X"E8",X"88",X"E8",
		X"02",X"27",X"E8",X"10",X"E8",X"02",X"EF",X"F8",X"10",X"F8",X"AA",X"00",X"7B",X"80",X"7B",X"A8",
		X"00",X"7B",X"D0",X"7B",X"F8",X"00",X"33",X"58",X"33",X"80",X"00",X"53",X"58",X"53",X"80",X"00",
		X"AB",X"58",X"AB",X"80",X"00",X"CB",X"58",X"CB",X"80",X"00",X"2B",X"80",X"2B",X"A8",X"00",X"D3",
		X"80",X"D3",X"A8",X"00",X"23",X"A8",X"23",X"D0",X"00",X"5B",X"A8",X"5B",X"D0",X"00",X"A3",X"A8",
		X"A3",X"D0",X"00",X"DB",X"A8",X"DB",X"D0",X"00",X"1B",X"D0",X"1B",X"F8",X"00",X"E3",X"D0",X"E3",
		X"F8",X"05",X"B7",X"30",X"48",X"30",X"05",X"CF",X"58",X"30",X"58",X"05",X"D7",X"80",X"28",X"80",
		X"05",X"DF",X"A8",X"20",X"A8",X"05",X"E7",X"D0",X"18",X"D0",X"05",X"EF",X"F8",X"10",X"F8",X"AA",
		X"FD",X"02",X"05",X"1D",X"FD",X"05",X"00",X"1D",X"FD",X"07",X"05",X"1D",X"01",X"00",X"00",X"1D",
		X"01",X"02",X"05",X"1D",X"01",X"05",X"00",X"1D",X"05",X"88",X"93",X"01",X"68",X"93",X"01",X"6C",
		X"93",X"03",X"49",X"93",X"05",X"08",X"93",X"01",X"E8",X"92",X"01",X"EC",X"92",X"05",X"C8",X"92",
		X"05",X"88",X"92",X"02",X"69",X"92",X"02",X"4A",X"92",X"05",X"28",X"92",X"05",X"E8",X"91",X"01",
		X"CA",X"91",X"03",X"A9",X"91",X"01",X"88",X"91",X"01",X"8C",X"91",X"05",X"48",X"91",X"01",X"28",
		X"91",X"01",X"2A",X"91",X"01",X"2C",X"91",X"01",X"08",X"91",X"01",X"0A",X"91",X"01",X"0C",X"91",
		X"03",X"C8",X"90",X"03",X"AA",X"90",X"03",X"88",X"90",X"05",X"2F",X"93",X"05",X"0F",X"93",X"02",
		X"F0",X"92",X"02",X"CF",X"92",X"02",X"D2",X"92",X"05",X"8F",X"92",X"05",X"6F",X"92",X"01",X"4F",
		X"92",X"01",X"53",X"92",X"05",X"2F",X"92",X"05",X"EF",X"91",X"02",X"D0",X"91",X"02",X"B1",X"91",
		X"05",X"8F",X"91",X"03",X"50",X"91",X"05",X"2F",X"91",X"01",X"0F",X"91",X"01",X"13",X"91",X"01",
		X"EF",X"90",X"01",X"F1",X"90",X"01",X"F3",X"90",X"02",X"D1",X"90",X"00",X"00",X"00",X"23",X"68",
		X"01",X"11",X"00",X"00",X"00",X"10",X"DB",X"68",X"01",X"40",X"00",X"00",X"08",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"01",X"C0",X"FF",
		X"01",X"FF",X"FF",X"34",X"C3",X"39",X"00",X"67",X"80",X"69",X"1A",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"04",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"1E",X"18",X"0B",X"4B",
		X"14",X"18",X"0B",X"4B",X"1E",X"18",X"0B",X"3B",X"14",X"18",X"0B",X"3B",X"3D",X"01",X"03",X"02",
		X"3D",X"01",X"04",X"01",X"27",X"70",X"01",X"E0",X"00",X"00",X"7F",X"40",X"01",X"78",X"02",X"00",
		X"27",X"49",X"0C",X"F0",X"7F",X"49",X"0C",X"88",X"1E",X"18",X"03",X"09",X"24",X"64",X"BB",X"C0",
		X"23",X"8D",X"7B",X"B4",X"1B",X"8C",X"7C",X"64",X"25",X"0E",X"04",X"02",X"23",X"46",X"03",X"68",
		X"DB",X"46",X"03",X"68",X"17",X"50",X"00",X"5C",X"E7",X"D0",X"00",X"5C",X"8C",X"50",X"00",X"84",
		X"73",X"D0",X"00",X"84",X"17",X"50",X"00",X"D4",X"E7",X"D0",X"00",X"D4",X"53",X"73",X"0A",X"A0",
		X"8B",X"74",X"0A",X"F0",X"DB",X"75",X"0A",X"A0",X"5B",X"73",X"0A",X"C8",X"E3",X"74",X"0A",X"60",
		X"1B",X"75",X"0A",X"80",X"DB",X"73",X"0A",X"C8",X"93",X"74",X"0A",X"F0",X"33",X"75",X"0A",X"50",
		X"1F",X"28",X"08",X"04",X"37",X"F4",X"37",X"C0",X"37",X"8C",X"77",X"70",X"77",X"A4",X"77",X"D8",
		X"11",X"01",X"00",X"06",X"2F",X"1F",X"D2",X"28",X"1E",X"1E",X"03",X"06",X"33",X"1F",X"D2",X"28",
		X"1E",X"1E",X"05",X"06",X"7F",X"C3",X"28",X"1E",X"3A",X"27",X"62",X"E5",X"EF",X"00",X"00",X"99",
		X"3E",X"B0",X"28",X"E0",X"28",X"01",X"29",X"00",X"00",X"E1",X"AF",X"32",X"60",X"60",X"06",X"04",
		X"11",X"20",X"00",X"DD",X"21",X"00",X"67",X"CD",X"C3",X"3E",X"00",X"00",X"CD",X"DC",X"42",X"00",
		X"CD",X"C3",X"3E",X"3A",X"60",X"60",X"A7",X"C8",X"FE",X"01",X"C8",X"FE",X"03",X"3E",X"03",X"D8",
		X"3E",X"07",X"C9",X"DD",X"CB",X"00",X"46",X"CA",X"FA",X"3E",X"79",X"DD",X"96",X"05",X"D2",X"D3",
		X"3E",X"ED",X"44",X"3C",X"95",X"DA",X"DE",X"3E",X"DD",X"96",X"0A",X"D2",X"FA",X"3E",X"FD",X"7E",
		X"03",X"DD",X"96",X"03",X"D2",X"E9",X"3E",X"ED",X"44",X"94",X"DA",X"F3",X"3E",X"DD",X"96",X"09",
		X"D2",X"FA",X"3E",X"3A",X"60",X"60",X"3C",X"32",X"60",X"60",X"DD",X"19",X"10",X"C5",X"C9",X"00",
		X"06",X"08",X"7E",X"12",X"23",X"13",X"7E",X"12",X"23",X"13",X"7E",X"D6",X"08",X"12",X"23",X"13",
		X"7E",X"D6",X"08",X"12",X"23",X"13",X"05",X"C2",X"02",X"3F",X"C9",X"21",X"C0",X"60",X"06",X"40",
		X"3E",X"FF",X"77",X"23",X"10",X"FC",X"21",X"00",X"88",X"06",X"00",X"77",X"23",X"10",X"FC",X"C3",
		X"9C",X"02",X"11",X"70",X"69",X"01",X"20",X"00",X"ED",X"B0",X"C9",X"DD",X"86",X"0F",X"77",X"CD",
		X"C0",X"46",X"C9",X"23",X"10",X"24",X"01",X"2C",X"6A",X"36",X"39",X"E5",X"2C",X"2C",X"7E",X"E1",
		X"C9",X"21",X"5D",X"93",X"3E",X"10",X"77",X"2C",X"77",X"01",X"20",X"00",X"09",X"77",X"2B",X"77",
		X"C9",X"FE",X"68",X"E1",X"CC",X"2E",X"3F",X"05",X"C2",X"15",X"29",X"AF",X"DD",X"E1",X"C9",X"3E",
		X"0A",X"90",X"FE",X"06",X"D8",X"C3",X"C5",X"2C",X"E6",X"F8",X"47",X"07",X"E6",X"10",X"4F",X"78",
		X"0F",X"0F",X"E6",X"04",X"B1",X"4F",X"78",X"0F",X"0F",X"E6",X"08",X"B1",X"4F",X"78",X"07",X"07",
		X"07",X"E6",X"02",X"B1",X"4F",X"78",X"07",X"E6",X"01",X"B1",X"C9",X"00",X"4C",X"49",X"4D",X"2E",
		X"CD",X"A6",X"3F",X"C3",X"5F",X"0D",X"3E",X"02",X"F7",X"06",X"02",X"21",X"6C",X"93",X"36",X"10",
		X"23",X"23",X"36",X"C0",X"21",X"8C",X"90",X"10",X"F5",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"7D",X"69",X"36",X"03",X"2C",X"2C",X"C9",X"06",X"08",X"21",X"00",X"60",X"AF",X"4F",X"77",
		X"23",X"0D",X"20",X"FB",X"10",X"F8",X"06",X"04",X"21",X"00",X"68",X"4F",X"77",X"23",X"0D",X"20",
		X"FB",X"10",X"F8",X"C3",X"74",X"02",X"0D",X"C2",X"67",X"0F",X"0E",X"03",X"16",X"00",X"21",X"00",
		X"68",X"42",X"77",X"23",X"10",X"FC",X"0D",X"20",X"F8",X"C3",X"6F",X"0F",X"7F",X"41",X"00",X"00",
		X"3A",X"27",X"62",X"C3",X"49",X"46",X"21",X"02",X"92",X"C3",X"E9",X"45",X"21",X"02",X"92",X"CD",
		X"A4",X"41",X"21",X"07",X"92",X"CD",X"E9",X"45",X"CD",X"35",X"40",X"C9",X"89",X"42",X"C9",X"32",
		X"00",X"93",X"21",X"80",X"9C",X"01",X"20",X"00",X"16",X"1A",X"3E",X"0C",X"CD",X"4E",X"40",X"21",
		X"81",X"9C",X"C3",X"46",X"40",X"21",X"42",X"91",X"3E",X"A0",X"CD",X"78",X"42",X"21",X"42",X"9D",
		X"3E",X"01",X"CD",X"89",X"42",X"C9",X"16",X"1A",X"3E",X"00",X"C3",X"B8",X"46",X"C9",X"77",X"09",
		X"15",X"20",X"FB",X"C9",X"21",X"42",X"91",X"3E",X"A4",X"CD",X"78",X"42",X"3E",X"01",X"21",X"42",
		X"9D",X"CD",X"89",X"42",X"C9",X"3A",X"26",X"60",X"A7",X"C0",X"21",X"DF",X"98",X"C3",X"A7",X"48",
		X"2B",X"77",X"C9",X"21",X"5D",X"93",X"3E",X"B4",X"CD",X"78",X"42",X"21",X"5D",X"9F",X"3E",X"0F",
		X"CD",X"89",X"42",X"C9",X"3E",X"0F",X"21",X"5D",X"9F",X"00",X"77",X"2C",X"77",X"09",X"77",X"2B",
		X"77",X"C9",X"21",X"46",X"93",X"CD",X"C3",X"40",X"21",X"48",X"93",X"CD",X"C3",X"40",X"21",X"86",
		X"93",X"CD",X"C3",X"40",X"21",X"88",X"93",X"CD",X"C3",X"40",X"21",X"46",X"9F",X"CD",X"C9",X"40",
		X"21",X"48",X"9F",X"CD",X"C9",X"40",X"21",X"86",X"9F",X"CD",X"C9",X"40",X"21",X"88",X"9F",X"CD",
		X"C9",X"40",X"C9",X"3E",X"60",X"CD",X"78",X"42",X"C9",X"3E",X"18",X"CD",X"89",X"42",X"C9",X"11",
		X"20",X"00",X"06",X"1E",X"21",X"48",X"9C",X"CD",X"F5",X"47",X"21",X"23",X"9D",X"06",X"16",X"CD",
		X"05",X"48",X"C3",X"CA",X"59",X"3A",X"26",X"60",X"A7",X"C0",X"21",X"DF",X"98",X"C3",X"84",X"48",
		X"C9",X"21",X"03",X"9E",X"3E",X"00",X"06",X"04",X"77",X"2C",X"10",X"FC",X"01",X"20",X"00",X"09",
		X"06",X"04",X"00",X"2B",X"10",X"FC",X"3A",X"00",X"62",X"C9",X"CD",X"F1",X"40",X"C9",X"03",X"92",
		X"E5",X"3E",X"FD",X"CD",X"89",X"42",X"E1",X"23",X"23",X"CD",X"89",X"42",X"C9",X"04",X"77",X"2B",
		X"10",X"FC",X"C9",X"21",X"46",X"93",X"3E",X"FD",X"C9",X"89",X"42",X"21",X"48",X"93",X"CD",X"89",
		X"42",X"21",X"86",X"93",X"CD",X"89",X"42",X"21",X"88",X"93",X"CD",X"89",X"42",X"C9",X"3E",X"B0",
		X"32",X"0C",X"92",X"32",X"2C",X"92",X"32",X"1E",X"92",X"32",X"3E",X"92",X"32",X"1E",X"93",X"32",
		X"3E",X"93",X"32",X"0C",X"93",X"32",X"2C",X"93",X"11",X"0F",X"00",X"C9",X"CA",X"06",X"40",X"21",
		X"03",X"92",X"C3",X"E9",X"45",X"CD",X"F0",X"45",X"CD",X"D6",X"46",X"21",X"90",X"63",X"C9",X"49",
		X"C3",X"F0",X"49",X"CD",X"23",X"41",X"CD",X"F1",X"40",X"C9",X"32",X"8B",X"63",X"CD",X"23",X"41",
		X"CD",X"F0",X"41",X"C9",X"CB",X"68",X"C2",X"8D",X"41",X"CD",X"77",X"48",X"C9",X"CD",X"8D",X"48",
		X"C9",X"23",X"36",X"F5",X"09",X"36",X"F7",X"2B",X"36",X"F6",X"01",X"E0",X"0B",X"09",X"3E",X"10",
		X"CD",X"89",X"42",X"C9",X"CD",X"10",X"41",X"21",X"02",X"9E",X"CD",X"F4",X"40",X"C9",X"21",X"5B",
		X"93",X"36",X"F8",X"23",X"36",X"F9",X"09",X"36",X"FB",X"2B",X"36",X"FA",X"01",X"E0",X"0B",X"09",
		X"3E",X"10",X"CD",X"89",X"42",X"C9",X"20",X"00",X"09",X"77",X"2B",X"77",X"00",X"00",X"00",X"C9",
		X"21",X"5B",X"93",X"01",X"20",X"00",X"3E",X"10",X"77",X"23",X"77",X"09",X"77",X"2B",X"77",X"01",
		X"E0",X"0B",X"09",X"3E",X"00",X"77",X"23",X"77",X"01",X"20",X"00",X"09",X"77",X"2B",X"77",X"C9",
		X"CD",X"0A",X"41",X"CD",X"D0",X"41",X"C9",X"21",X"DF",X"98",X"36",X"13",X"2B",X"36",X"00",X"2B",
		X"36",X"12",X"21",X"55",X"88",X"36",X"FF",X"2C",X"36",X"FF",X"2C",X"36",X"30",X"2C",X"36",X"31",
		X"01",X"10",X"00",X"09",X"36",X"33",X"2B",X"36",X"32",X"2B",X"36",X"FF",X"2B",X"36",X"FF",X"09",
		X"36",X"3C",X"2C",X"36",X"3D",X"2C",X"36",X"38",X"2C",X"36",X"39",X"09",X"36",X"3B",X"2B",X"36",
		X"3A",X"2B",X"36",X"3F",X"2B",X"36",X"3E",X"09",X"36",X"40",X"2C",X"36",X"41",X"2C",X"36",X"34",
		X"2C",X"36",X"35",X"09",X"36",X"37",X"2B",X"36",X"36",X"2B",X"36",X"43",X"2B",X"36",X"42",X"C9",
		X"21",X"DD",X"98",X"36",X"22",X"C9",X"21",X"18",X"91",X"3E",X"78",X"CD",X"78",X"42",X"21",X"18",
		X"9D",X"3E",X"10",X"CD",X"89",X"42",X"00",X"21",X"6C",X"93",X"3E",X"78",X"CD",X"78",X"42",X"21",
		X"6C",X"9F",X"3E",X"10",X"CD",X"89",X"42",X"C9",X"C5",X"77",X"2C",X"3C",X"77",X"01",X"20",X"00",
		X"09",X"3C",X"3C",X"77",X"2B",X"3D",X"77",X"C1",X"C9",X"C5",X"77",X"2C",X"77",X"01",X"20",X"00",
		X"09",X"77",X"2B",X"77",X"C1",X"C9",X"00",X"00",X"00",X"3A",X"81",X"66",X"E6",X"01",X"C2",X"B2",
		X"42",X"21",X"18",X"91",X"3E",X"FD",X"CD",X"89",X"42",X"21",X"18",X"9D",X"3E",X"00",X"CD",X"89",
		X"42",X"C9",X"21",X"6C",X"93",X"3E",X"FD",X"CD",X"89",X"42",X"21",X"6C",X"9F",X"3E",X"00",X"CD",
		X"89",X"42",X"C9",X"11",X"78",X"69",X"3A",X"27",X"62",X"FE",X"01",X"C2",X"D1",X"42",X"06",X"01",
		X"C9",X"FE",X"04",X"C2",X"75",X"45",X"06",X"05",X"C9",X"06",X"02",X"C9",X"DD",X"21",X"00",X"64",
		X"C3",X"C6",X"42",X"11",X"20",X"00",X"C3",X"C6",X"42",X"CD",X"C6",X"42",X"78",X"C9",X"3E",X"06",
		X"90",X"D8",X"C3",X"DC",X"25",X"3E",X"07",X"85",X"6F",X"C9",X"3A",X"27",X"62",X"FE",X"01",X"CA",
		X"56",X"42",X"FE",X"02",X"CA",X"28",X"43",X"21",X"EC",X"91",X"3E",X"78",X"CD",X"78",X"42",X"21",
		X"EC",X"9D",X"3E",X"10",X"CD",X"89",X"42",X"21",X"71",X"93",X"3E",X"14",X"CD",X"78",X"42",X"21",
		X"71",X"9F",X"3E",X"20",X"CD",X"89",X"42",X"C9",X"21",X"F6",X"91",X"3E",X"78",X"CD",X"78",X"42",
		X"21",X"F6",X"9D",X"3E",X"10",X"CD",X"89",X"42",X"21",X"71",X"93",X"3E",X"14",X"CD",X"78",X"42",
		X"21",X"71",X"9F",X"3E",X"20",X"CD",X"89",X"42",X"C9",X"E5",X"F5",X"D6",X"68",X"07",X"21",X"7F",
		X"43",X"06",X"00",X"4F",X"09",X"F1",X"C2",X"6C",X"43",X"7E",X"32",X"6D",X"93",X"23",X"7E",X"32",
		X"6C",X"93",X"3E",X"24",X"32",X"6C",X"9F",X"32",X"6D",X"9F",X"E1",X"C9",X"7E",X"32",X"8D",X"90",
		X"23",X"7E",X"32",X"8C",X"90",X"3E",X"24",X"32",X"8C",X"9C",X"32",X"8D",X"9C",X"E1",X"C9",X"1F",
		X"1F",X"1F",X"1E",X"1F",X"1D",X"1F",X"1C",X"1F",X"1B",X"1F",X"1A",X"1F",X"19",X"1F",X"18",X"1F",
		X"FD",X"1F",X"FD",X"1E",X"FD",X"1D",X"FD",X"1C",X"FD",X"1B",X"FD",X"1A",X"FD",X"19",X"FD",X"FD",
		X"FD",X"21",X"93",X"92",X"3E",X"94",X"CD",X"78",X"42",X"21",X"93",X"9E",X"3E",X"01",X"CD",X"89",
		X"42",X"21",X"73",X"90",X"3E",X"9C",X"CD",X"78",X"42",X"21",X"73",X"9C",X"3E",X"01",X"CD",X"89",
		X"42",X"21",X"FD",X"91",X"3E",X"98",X"CD",X"78",X"42",X"21",X"FD",X"9D",X"3E",X"01",X"CD",X"89",
		X"42",X"21",X"F0",X"91",X"3E",X"B4",X"CD",X"78",X"42",X"21",X"F0",X"9D",X"3E",X"02",X"CD",X"89",
		X"42",X"C9",X"21",X"8F",X"93",X"3E",X"9C",X"CD",X"78",X"42",X"21",X"8F",X"9F",X"3E",X"01",X"CD",
		X"89",X"42",X"21",X"4B",X"90",X"3E",X"98",X"CD",X"78",X"42",X"21",X"4B",X"9C",X"3E",X"01",X"CD",
		X"89",X"42",X"21",X"98",X"92",X"3E",X"4C",X"CD",X"78",X"42",X"21",X"98",X"9E",X"3E",X"04",X"CD",
		X"89",X"42",X"C9",X"21",X"09",X"93",X"3E",X"9C",X"CD",X"78",X"42",X"21",X"09",X"9F",X"3E",X"01",
		X"CD",X"89",X"42",X"21",X"7D",X"91",X"3E",X"98",X"CD",X"78",X"42",X"21",X"7D",X"9D",X"3E",X"01",
		X"CD",X"89",X"42",X"21",X"78",X"90",X"3E",X"4C",X"CD",X"78",X"42",X"21",X"78",X"9C",X"3E",X"04",
		X"CD",X"89",X"42",X"C9",X"3E",X"11",X"32",X"07",X"9E",X"21",X"25",X"6A",X"C9",X"CD",X"C0",X"47",
		X"C3",X"95",X"13",X"20",X"00",X"09",X"36",X"47",X"2B",X"36",X"46",X"2B",X"36",X"43",X"2B",X"36",
		X"42",X"21",X"07",X"9E",X"3E",X"10",X"CD",X"89",X"42",X"21",X"0A",X"9E",X"C3",X"68",X"46",X"C9",
		X"3E",X"FD",X"CD",X"89",X"42",X"C3",X"E0",X"59",X"09",X"3E",X"00",X"CD",X"89",X"42",X"C9",X"36",
		X"FD",X"23",X"36",X"10",X"01",X"20",X"00",X"09",X"36",X"C0",X"2B",X"36",X"C0",X"C9",X"00",X"00",
		X"21",X"02",X"92",X"CD",X"70",X"44",X"21",X"04",X"92",X"C3",X"70",X"44",X"21",X"73",X"90",X"C3",
		X"70",X"44",X"21",X"FD",X"91",X"C3",X"70",X"44",X"21",X"93",X"92",X"C3",X"70",X"44",X"21",X"F0",
		X"91",X"C3",X"70",X"44",X"21",X"8F",X"93",X"C3",X"70",X"44",X"21",X"4B",X"90",X"C3",X"70",X"44",
		X"21",X"98",X"92",X"C3",X"EB",X"59",X"21",X"09",X"93",X"C3",X"70",X"44",X"21",X"7D",X"91",X"C3",
		X"70",X"44",X"21",X"78",X"90",X"C3",X"EB",X"59",X"32",X"B9",X"62",X"CD",X"A1",X"43",X"C9",X"DD",
		X"21",X"00",X"64",X"CD",X"E2",X"43",X"C9",X"11",X"A3",X"64",X"CD",X"13",X"44",X"C9",X"22",X"43",
		X"63",X"7D",X"FE",X"0C",X"CA",X"1C",X"45",X"FE",X"10",X"CA",X"0C",X"45",X"3A",X"27",X"62",X"FE",
		X"02",X"CA",X"9C",X"44",X"FE",X"03",X"CA",X"B4",X"44",X"C3",X"C6",X"44",X"3A",X"27",X"62",X"FE",
		X"02",X"CA",X"A2",X"44",X"FE",X"03",X"CA",X"BA",X"44",X"C3",X"CC",X"44",X"3A",X"27",X"62",X"FE",
		X"02",X"CA",X"A8",X"44",X"FE",X"03",X"CA",X"C0",X"44",X"C3",X"D2",X"44",X"3E",X"2B",X"32",X"4B",
		X"9C",X"32",X"5A",X"9C",X"32",X"D0",X"9D",X"32",X"30",X"9E",X"32",X"AB",X"9F",X"32",X"BA",X"9F",
		X"2C",X"1A",X"17",X"C9",X"FE",X"AB",X"C2",X"4D",X"45",X"21",X"4B",X"90",X"C9",X"FE",X"D0",X"C2",
		X"56",X"45",X"21",X"30",X"92",X"C9",X"21",X"5A",X"90",X"C9",X"CD",X"2C",X"45",X"3E",X"21",X"32",
		X"4B",X"90",X"32",X"5A",X"90",X"32",X"D0",X"91",X"32",X"30",X"92",X"32",X"AB",X"93",X"32",X"BA",
		X"93",X"21",X"18",X"3E",X"C9",X"FE",X"03",X"C2",X"52",X"01",X"06",X"01",X"C9",X"E5",X"23",X"23",
		X"77",X"E1",X"C3",X"BB",X"25",X"CD",X"F0",X"45",X"DF",X"0E",X"17",X"C3",X"92",X"13",X"41",X"41",
		X"21",X"55",X"88",X"3E",X"80",X"CD",X"47",X"49",X"3E",X"8C",X"CD",X"47",X"49",X"3E",X"98",X"CD",
		X"47",X"49",X"21",X"57",X"88",X"3E",X"84",X"CD",X"47",X"49",X"3E",X"90",X"CD",X"47",X"49",X"3E",
		X"9C",X"CD",X"47",X"49",X"21",X"59",X"88",X"3E",X"88",X"CD",X"47",X"49",X"3E",X"94",X"CD",X"47",
		X"49",X"3E",X"A0",X"CD",X"47",X"49",X"3E",X"01",X"32",X"00",X"6B",X"C9",X"A7",X"7E",X"ED",X"52",
		X"FE",X"19",X"D2",X"DB",X"45",X"23",X"23",X"36",X"00",X"2B",X"2B",X"2B",X"05",X"C8",X"C3",X"CC",
		X"45",X"CD",X"6C",X"17",X"13",X"23",X"23",X"23",X"C9",X"E5",X"E5",X"C3",X"E2",X"4F",X"41",X"41",
		X"21",X"00",X"88",X"06",X"00",X"3E",X"FF",X"77",X"23",X"10",X"FC",X"C9",X"CD",X"89",X"42",X"C9",
		X"E5",X"CD",X"78",X"42",X"01",X"00",X"0C",X"E1",X"09",X"3E",X"2B",X"CD",X"89",X"42",X"C9",X"41",
		X"C3",X"60",X"47",X"FE",X"01",X"20",X"09",X"21",X"5B",X"93",X"3E",X"00",X"CD",X"00",X"46",X"C9",
		X"21",X"EE",X"91",X"3E",X"00",X"C3",X"54",X"47",X"C9",X"21",X"DD",X"98",X"C3",X"B9",X"47",X"3B",
		X"C3",X"74",X"47",X"FE",X"01",X"20",X"09",X"21",X"5B",X"93",X"3E",X"08",X"CD",X"00",X"46",X"C9",
		X"21",X"EE",X"91",X"3E",X"08",X"C3",X"54",X"47",X"C9",X"FE",X"04",X"C3",X"5C",X"41",X"41",X"41",
		X"36",X"4D",X"23",X"36",X"4C",X"01",X"20",X"00",X"09",X"36",X"4E",X"2C",X"36",X"4F",X"01",X"E0",
		X"0B",X"09",X"3E",X"20",X"CD",X"89",X"42",X"C9",X"CD",X"89",X"42",X"C3",X"77",X"46",X"41",X"41",
		X"CD",X"74",X"08",X"CD",X"F0",X"45",X"C9",X"CD",X"0A",X"41",X"CD",X"35",X"40",X"C9",X"2B",X"41",
		X"CD",X"A3",X"49",X"3A",X"10",X"69",X"C9",X"CD",X"F0",X"45",X"DF",X"0E",X"17",X"C3",X"A4",X"13",
		X"C5",X"CB",X"68",X"C2",X"A8",X"46",X"CD",X"10",X"46",X"3A",X"27",X"62",X"C1",X"FE",X"01",X"CA",
		X"84",X"41",X"CD",X"C2",X"48",X"C9",X"00",X"00",X"CD",X"30",X"46",X"3A",X"27",X"62",X"FE",X"01",
		X"C1",X"CA",X"84",X"41",X"CD",X"B5",X"48",X"C9",X"CD",X"4E",X"40",X"CD",X"C0",X"47",X"C9",X"41",
		X"DD",X"77",X"05",X"3A",X"27",X"62",X"FE",X"01",X"CA",X"99",X"42",X"FE",X"02",X"28",X"29",X"3A",
		X"81",X"66",X"E6",X"01",X"20",X"11",X"21",X"EC",X"91",X"3E",X"FD",X"CD",X"89",X"42",X"21",X"EC",
		X"9D",X"3E",X"00",X"CD",X"89",X"42",X"C9",X"21",X"71",X"93",X"3E",X"FD",X"CD",X"89",X"42",X"21",
		X"71",X"9F",X"3E",X"00",X"CD",X"89",X"42",X"C9",X"3A",X"81",X"66",X"E6",X"01",X"20",X"11",X"21",
		X"F6",X"91",X"3E",X"FD",X"CD",X"89",X"42",X"21",X"F6",X"9D",X"3E",X"00",X"CD",X"89",X"42",X"C9",
		X"21",X"71",X"93",X"3E",X"FD",X"CD",X"89",X"42",X"3E",X"00",X"21",X"71",X"9F",X"CD",X"89",X"42",
		X"C9",X"CD",X"9A",X"48",X"21",X"EC",X"3D",X"C9",X"3A",X"27",X"62",X"FE",X"02",X"C0",X"C3",X"80",
		X"46",X"3A",X"27",X"62",X"FE",X"04",X"C2",X"90",X"46",X"3E",X"40",X"32",X"DE",X"98",X"C3",X"90",
		X"46",X"CD",X"86",X"11",X"CD",X"21",X"47",X"C9",X"CD",X"21",X"47",X"3E",X"40",X"32",X"DE",X"98",
		X"21",X"F0",X"3D",X"C9",X"C3",X"00",X"46",X"21",X"5B",X"93",X"3E",X"FD",X"CD",X"89",X"42",X"C9",
		X"3A",X"27",X"62",X"FE",X"04",X"C8",X"FE",X"03",X"C2",X"13",X"46",X"21",X"EE",X"91",X"3E",X"FD",
		X"CD",X"89",X"42",X"C9",X"3A",X"27",X"62",X"FE",X"04",X"C8",X"FE",X"03",X"C2",X"33",X"46",X"C3",
		X"6B",X"47",X"23",X"41",X"41",X"DD",X"2A",X"51",X"63",X"16",X"00",X"3A",X"53",X"63",X"5F",X"01",
		X"04",X"00",X"3A",X"54",X"63",X"A7",X"CA",X"A0",X"47",X"09",X"DD",X"19",X"3D",X"C2",X"99",X"47",
		X"DD",X"36",X"00",X"00",X"DD",X"7E",X"15",X"A7",X"3E",X"02",X"CA",X"AF",X"47",X"3E",X"04",X"32",
		X"42",X"63",X"23",X"36",X"1E",X"2B",X"C3",X"E1",X"1E",X"36",X"BB",X"23",X"C3",X"F0",X"47",X"25",
		X"F5",X"C5",X"D5",X"E5",X"3A",X"27",X"62",X"FE",X"01",X"20",X"06",X"3E",X"0A",X"C3",X"CF",X"40",
		X"C9",X"FE",X"02",X"20",X"06",X"3E",X"04",X"C3",X"CF",X"40",X"C9",X"FE",X"03",X"20",X"06",X"3E",
		X"06",X"C3",X"CF",X"40",X"C9",X"3E",X"02",X"C3",X"CF",X"40",X"00",X"E1",X"D1",X"C1",X"F1",X"C9",
		X"36",X"98",X"C3",X"1C",X"48",X"0E",X"18",X"E5",X"77",X"0D",X"23",X"20",X"FB",X"E1",X"19",X"10",
		X"F4",X"C9",X"2D",X"41",X"41",X"0E",X"06",X"E5",X"77",X"0D",X"23",X"20",X"FB",X"E1",X"19",X"10",
		X"F4",X"C9",X"CD",X"70",X"48",X"CD",X"F0",X"45",X"21",X"09",X"60",X"C9",X"23",X"36",X"A0",X"C9",
		X"CD",X"C0",X"47",X"3A",X"27",X"62",X"C9",X"41",X"41",X"3F",X"CD",X"2A",X"12",X"CD",X"C0",X"47",
		X"C9",X"41",X"CD",X"32",X"3F",X"C9",X"D6",X"46",X"C3",X"E5",X"48",X"E5",X"48",X"CD",X"C0",X"47",
		X"21",X"F0",X"3C",X"C9",X"41",X"CD",X"77",X"48",X"11",X"07",X"68",X"C9",X"2B",X"41",X"41",X"41",
		X"D5",X"32",X"01",X"A0",X"32",X"02",X"A0",X"36",X"03",X"32",X"01",X"6B",X"D1",X"C9",X"41",X"41",
		X"32",X"01",X"A0",X"32",X"02",X"A0",X"32",X"01",X"6B",X"C9",X"CD",X"C0",X"47",X"C3",X"D5",X"48",
		X"CD",X"C0",X"47",X"CD",X"16",X"06",X"C9",X"3A",X"01",X"6B",X"A7",X"C2",X"F7",X"41",X"CD",X"F7",
		X"41",X"C3",X"E5",X"40",X"36",X"7B",X"2B",X"36",X"00",X"2B",X"36",X"02",X"C9",X"3A",X"01",X"6B",
		X"A7",X"C3",X"E2",X"07",X"21",X"DD",X"98",X"36",X"32",X"C9",X"3A",X"01",X"6B",X"A7",X"C2",X"58",
		X"49",X"CD",X"58",X"49",X"C3",X"65",X"40",X"36",X"80",X"2B",X"36",X"01",X"2B",X"36",X"02",X"3E",
		X"00",X"32",X"00",X"6B",X"C9",X"3A",X"26",X"60",X"A7",X"C3",X"BB",X"4F",X"21",X"DD",X"98",X"36",
		X"32",X"C9",X"3A",X"26",X"60",X"A7",X"C3",X"C8",X"4F",X"21",X"DD",X"98",X"36",X"12",X"C9",X"32",
		X"01",X"6B",X"36",X"03",X"C9",X"21",X"00",X"69",X"C9",X"41",X"06",X"02",X"77",X"19",X"00",X"10",
		X"FB",X"C9",X"41",X"39",X"29",X"CD",X"C0",X"47",X"11",X"CF",X"39",X"C9",X"41",X"41",X"CD",X"C0",
		X"47",X"21",X"48",X"60",X"C9",X"CD",X"C9",X"45",X"CD",X"F0",X"45",X"C9",X"CD",X"F0",X"45",X"DF",
		X"D5",X"06",X"11",X"2A",X"E4",X"69",X"11",X"11",X"00",X"19",X"22",X"E4",X"69",X"11",X"FA",X"48",
		X"ED",X"52",X"7C",X"E6",X"80",X"CA",X"25",X"49",X"2A",X"E4",X"69",X"D1",X"7E",X"CD",X"E2",X"49",
		X"50",X"C2",X"1C",X"49",X"C9",X"21",X"75",X"45",X"22",X"E4",X"69",X"C3",X"1C",X"49",X"11",X"0D",
		X"93",X"21",X"75",X"45",X"22",X"E4",X"69",X"CD",X"00",X"49",X"21",X"0D",X"9F",X"06",X"11",X"36",
		X"20",X"23",X"05",X"C2",X"3F",X"49",X"C9",X"C5",X"77",X"23",X"3C",X"77",X"01",X"10",X"00",X"09",
		X"3C",X"3C",X"77",X"3D",X"2B",X"C3",X"6D",X"49",X"21",X"DF",X"98",X"36",X"10",X"2B",X"36",X"01",
		X"2B",X"36",X"12",X"C3",X"90",X"45",X"01",X"10",X"00",X"3E",X"88",X"D1",X"0A",X"77",X"09",X"C1",
		X"C9",X"3E",X"85",X"CD",X"47",X"49",X"3E",X"84",X"CD",X"47",X"49",X"3E",X"81",X"CD",X"47",X"49",
		X"3E",X"80",X"CD",X"47",X"49",X"ED",X"42",X"D1",X"05",X"00",X"19",X"36",X"FF",X"ED",X"42",X"36",
		X"FF",X"3E",X"00",X"32",X"00",X"6B",X"C9",X"21",X"DD",X"98",X"36",X"22",X"C9",X"21",X"DD",X"98",
		X"36",X"02",X"C9",X"21",X"DE",X"98",X"3A",X"00",X"6B",X"A7",X"28",X"0D",X"7E",X"3D",X"28",X"02",
		X"77",X"C9",X"3C",X"77",X"AF",X"32",X"00",X"6B",X"C9",X"7E",X"3C",X"FE",X"80",X"28",X"02",X"77",
		X"C9",X"3D",X"77",X"3E",X"01",X"32",X"00",X"6B",X"C9",X"F5",X"E5",X"21",X"01",X"A0",X"3E",X"01",
		X"77",X"23",X"77",X"3E",X"01",X"32",X"01",X"6B",X"E1",X"F1",X"C9",X"AF",X"77",X"23",X"77",X"E1",
		X"F1",X"C9",X"12",X"3C",X"E5",X"C5",X"01",X"20",X"00",X"EB",X"09",X"77",X"EB",X"C1",X"E1",X"C9",
		X"FE",X"03",X"CC",X"FC",X"49",X"ED",X"B0",X"C9",X"11",X"74",X"69",X"C9",X"11",X"7C",X"69",X"C9",
		X"21",X"FC",X"6B",X"3A",X"FF",X"6B",X"A7",X"20",X"20",X"21",X"89",X"60",X"CD",X"80",X"4E",X"00",
		X"00",X"00",X"00",X"7E",X"A7",X"20",X"06",X"21",X"88",X"60",X"C3",X"F0",X"4E",X"36",X"00",X"21",
		X"FE",X"6B",X"77",X"2D",X"AF",X"77",X"2D",X"3C",X"77",X"7E",X"3D",X"77",X"C0",X"2C",X"34",X"3A",
		X"FE",X"6B",X"21",X"E3",X"4A",X"87",X"CD",X"61",X"4A",X"5E",X"23",X"56",X"EB",X"22",X"FA",X"6B",
		X"3A",X"FD",X"6B",X"3D",X"C3",X"D0",X"4E",X"87",X"91",X"C6",X"06",X"CD",X"61",X"4A",X"7E",X"32",
		X"FF",X"6B",X"A7",X"C8",X"32",X"FC",X"6B",X"23",X"EB",X"2A",X"FA",X"6B",X"EB",X"CD",X"69",X"4A",
		X"C9",X"A7",X"85",X"6F",X"3E",X"00",X"8C",X"67",X"C9",X"00",X"00",X"00",X"CD",X"8D",X"4A",X"0E",
		X"00",X"CD",X"77",X"4A",X"EB",X"0E",X"08",X"06",X"06",X"79",X"D3",X"08",X"0C",X"7E",X"D3",X"09",
		X"23",X"10",X"F6",X"C9",X"3E",X"07",X"D3",X"08",X"3E",X"3F",X"D3",X"09",X"C9",X"3E",X"07",X"D3",
		X"08",X"3E",X"38",X"18",X"F5",X"87",X"21",X"D3",X"4A",X"CD",X"61",X"4A",X"7E",X"32",X"00",X"A8",
		X"AF",X"32",X"07",X"A0",X"3E",X"07",X"D3",X"08",X"3E",X"C0",X"D3",X"09",X"3E",X"0E",X"D3",X"08",
		X"23",X"7E",X"D3",X"09",X"3E",X"0F",X"D3",X"08",X"3E",X"7F",X"D3",X"09",X"3E",X"07",X"32",X"00",
		X"B0",X"32",X"04",X"A0",X"AF",X"32",X"04",X"A0",X"CD",X"70",X"4E",X"3E",X"FF",X"32",X"04",X"A0",
		X"C9",X"A0",X"C9",X"4F",X"40",X"79",X"28",X"70",X"C0",X"20",X"97",X"04",X"A5",X"7F",X"7F",X"C0",
		X"68",X"7C",X"70",X"03",X"4B",X"37",X"4C",X"61",X"4C",X"99",X"4C",X"A0",X"54",X"D1",X"4C",X"3A",
		X"4D",X"79",X"4D",X"E9",X"4D",X"F0",X"4D",X"F7",X"4D",X"FE",X"4D",X"8B",X"4E",X"0C",X"4E",X"36",
		X"4E",X"60",X"4E",X"1F",X"1F",X"1F",X"FF",X"0F",X"00",X"08",X"2D",X"00",X"2D",X"00",X"2D",X"00",
		X"10",X"2F",X"00",X"2F",X"00",X"2F",X"00",X"08",X"35",X"00",X"35",X"00",X"35",X"00",X"10",X"3C",
		X"00",X"3C",X"00",X"3C",X"00",X"08",X"43",X"00",X"43",X"00",X"43",X"00",X"10",X"47",X"00",X"47",
		X"00",X"47",X"00",X"08",X"50",X"00",X"50",X"00",X"50",X"00",X"10",X"5A",X"00",X"5A",X"00",X"5A",
		X"00",X"08",X"5F",X"00",X"5F",X"00",X"5F",X"00",X"10",X"6B",X"00",X"6B",X"00",X"6B",X"00",X"08",
		X"78",X"00",X"78",X"00",X"78",X"00",X"10",X"86",X"00",X"86",X"00",X"86",X"00",X"08",X"8E",X"00",
		X"8E",X"00",X"8E",X"00",X"10",X"A0",X"00",X"A0",X"00",X"A0",X"00",X"20",X"B3",X"00",X"B3",X"00",
		X"1C",X"01",X"10",X"B3",X"00",X"B3",X"00",X"3F",X"01",X"20",X"B3",X"00",X"B3",X"00",X"66",X"01",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"B6",X"4B",X"11",X"C2",X"92",X"0E",X"05",X"06",X"03",X"ED",X"B0",X"CD",X"C5",X"4B",X"0D",
		X"20",X"F6",X"11",X"C2",X"9E",X"3E",X"01",X"0E",X"05",X"06",X"03",X"12",X"13",X"10",X"FC",X"CD",
		X"C5",X"4B",X"0D",X"20",X"F4",X"C9",X"8A",X"FD",X"FD",X"87",X"88",X"89",X"84",X"85",X"86",X"81",
		X"82",X"83",X"80",X"FD",X"FD",X"E5",X"21",X"1C",X"00",X"19",X"EB",X"E1",X"C9",X"FF",X"FF",X"FF",
		X"21",X"D9",X"91",X"11",X"EE",X"4B",X"06",X"06",X"1A",X"77",X"E5",X"D5",X"11",X"00",X"0C",X"19",
		X"36",X"02",X"D1",X"E1",X"D5",X"11",X"20",X"00",X"19",X"D1",X"13",X"10",X"E8",X"C9",X"06",X"01",
		X"12",X"03",X"1F",X"1E",X"00",X"00",X"00",X"01",X"20",X"00",X"1E",X"05",X"16",X"0F",X"CD",X"07",
		X"4C",X"23",X"1D",X"C2",X"FC",X"4B",X"C9",X"E5",X"00",X"77",X"09",X"15",X"C2",X"09",X"4C",X"E1",
		X"C9",X"21",X"14",X"9D",X"3E",X"00",X"CD",X"F4",X"4B",X"3E",X"FD",X"21",X"14",X"91",X"CD",X"F4",
		X"4B",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"1F",X"FF",X"2F",X"00",X"60",X"66",X"01",
		X"5A",X"00",X"5A",X"00",X"1A",X"3F",X"01",X"50",X"00",X"50",X"00",X"38",X"2D",X"01",X"4B",X"00",
		X"2D",X"01",X"38",X"66",X"01",X"5A",X"00",X"5A",X"00",X"60",X"FD",X"00",X"40",X"00",X"EF",X"00",
		X"00",X"1F",X"1F",X"1F",X"87",X"17",X"00",X"20",X"B3",X"00",X"B3",X"00",X"B3",X"00",X"10",X"86",
		X"00",X"86",X"00",X"86",X"00",X"20",X"8E",X"00",X"8E",X"00",X"8E",X"00",X"10",X"78",X"00",X"78",
		X"00",X"78",X"00",X"10",X"86",X"00",X"86",X"00",X"86",X"00",X"10",X"6B",X"00",X"6B",X"00",X"6B",
		X"00",X"40",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"00",X"1F",X"1F",X"1F",X"98",X"0F",X"00",X"08",
		X"43",X"00",X"43",X"00",X"43",X"00",X"08",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"08",X"35",X"00",
		X"35",X"00",X"35",X"00",X"08",X"43",X"00",X"43",X"00",X"43",X"00",X"08",X"3C",X"00",X"3C",X"00",
		X"3C",X"00",X"08",X"35",X"00",X"35",X"00",X"35",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"00",
		X"00",X"1F",X"1F",X"1F",X"FF",X"22",X"00",X"20",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"20",X"2F",
		X"00",X"2F",X"00",X"2F",X"00",X"08",X"40",X"00",X"40",X"00",X"40",X"00",X"10",X"35",X"00",X"35",
		X"00",X"35",X"00",X"10",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"10",X"43",X"00",X"43",X"00",X"43",
		X"00",X"10",X"50",X"00",X"50",X"00",X"50",X"00",X"20",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"10",
		X"47",X"00",X"47",X"00",X"47",X"00",X"10",X"50",X"00",X"50",X"00",X"50",X"00",X"08",X"47",X"00",
		X"47",X"00",X"47",X"00",X"20",X"50",X"00",X"50",X"00",X"50",X"00",X"10",X"5A",X"00",X"5A",X"00",
		X"5A",X"00",X"80",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"00",X"1F",X"1F",X"1F",X"80",X"08",X"00",
		X"10",X"78",X"00",X"EF",X"00",X"78",X"00",X"04",X"6B",X"00",X"6B",X"00",X"6B",X"00",X"04",X"5F",
		X"00",X"5F",X"00",X"5F",X"00",X"04",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"04",X"50",X"00",X"50",
		X"00",X"50",X"00",X"04",X"47",X"00",X"47",X"00",X"47",X"00",X"04",X"43",X"00",X"43",X"00",X"43",
		X"00",X"04",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"00",X"1F",X"1F",X"1F",X"60",X"1A",X"00",X"08",
		X"6B",X"00",X"5F",X"00",X"6B",X"00",X"08",X"6B",X"00",X"5F",X"00",X"6B",X"00",X"10",X"6B",X"00",
		X"5F",X"00",X"6B",X"00",X"08",X"6B",X"00",X"5F",X"00",X"6B",X"00",X"08",X"5A",X"00",X"50",X"00",
		X"5A",X"00",X"08",X"5A",X"00",X"50",X"00",X"5A",X"00",X"10",X"5A",X"00",X"50",X"00",X"5A",X"00",
		X"08",X"5A",X"00",X"50",X"00",X"5A",X"00",X"08",X"47",X"00",X"43",X"00",X"47",X"00",X"08",X"47",
		X"00",X"43",X"00",X"47",X"00",X"10",X"47",X"00",X"43",X"00",X"47",X"00",X"08",X"47",X"00",X"43",
		X"00",X"47",X"00",X"10",X"66",X"01",X"66",X"01",X"66",X"01",X"10",X"1C",X"01",X"1C",X"01",X"1C",
		X"01",X"10",X"66",X"01",X"1C",X"01",X"EF",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"1F",X"1F",X"1F",X"40",
		X"11",X"00",X"04",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"04",X"50",X"00",X"50",X"00",X"50",X"00",
		X"04",X"47",X"00",X"47",X"00",X"47",X"00",X"04",X"43",X"00",X"43",X"00",X"43",X"00",X"04",X"3C",
		X"00",X"3C",X"00",X"3C",X"00",X"00",X"1F",X"1F",X"1F",X"33",X"1B",X"00",X"20",X"43",X"00",X"35",
		X"00",X"43",X"00",X"10",X"35",X"00",X"2D",X"00",X"35",X"00",X"10",X"35",X"00",X"2D",X"00",X"35",
		X"00",X"10",X"35",X"00",X"2D",X"00",X"35",X"00",X"20",X"35",X"00",X"2D",X"00",X"35",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"C5",X"01",X"80",X"02",X"0D",X"20",X"FD",X"10",X"FB",X"C1",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"8B",X"60",X"A7",X"C8",X"00",X"32",X"8B",X"60",X"2C",X"C9",X"1F",X"1F",X"1F",X"FF",X"4F",
		X"00",X"20",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"08",X"47",X"00",X"47",X"00",X"47",X"00",X"10",
		X"50",X"00",X"50",X"00",X"50",X"00",X"10",X"5A",X"00",X"5A",X"00",X"5A",X"00",X"10",X"43",X"00",
		X"43",X"00",X"43",X"00",X"10",X"3C",X"00",X"3C",X"00",X"3C",X"00",X"10",X"35",X"00",X"35",X"00",
		X"35",X"00",X"40",X"2F",X"00",X"2F",X"00",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EB",X"26",X"00",X"6F",X"29",X"29",X"29",X"D5",X"16",X"00",X"5F",X"A7",X"ED",X"52",X"1E",X"06",
		X"19",X"D1",X"19",X"C3",X"4E",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"A7",X"C8",X"AF",X"C3",X"1D",X"4A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"65",X"93",X"01",X"45",X"93",X"01",X"4A",X"93",X"01",X"25",X"93",X"01",X"2A",X"93",X"02",
		X"05",X"93",X"02",X"09",X"93",X"06",X"C6",X"92",X"01",X"A6",X"92",X"01",X"A9",X"92",X"01",X"86",
		X"92",X"02",X"89",X"92",X"04",X"66",X"92",X"01",X"6B",X"92",X"05",X"26",X"92",X"01",X"05",X"92",
		X"01",X"08",X"92",X"01",X"E5",X"91",X"01",X"E8",X"91",X"05",X"C6",X"91",X"01",X"86",X"91",X"02",
		X"8A",X"91",X"01",X"66",X"91",X"01",X"69",X"91",X"01",X"6B",X"91",X"01",X"46",X"91",X"01",X"48",
		X"91",X"01",X"4B",X"91",X"02",X"26",X"91",X"01",X"2B",X"91",X"03",X"E5",X"90",X"01",X"C8",X"90",
		X"03",X"A8",X"90",X"01",X"88",X"90",X"03",X"65",X"90",X"06",X"4E",X"93",X"06",X"2E",X"93",X"02",
		X"10",X"93",X"02",X"EE",X"92",X"02",X"F2",X"92",X"02",X"CE",X"92",X"02",X"D2",X"92",X"06",X"8E",
		X"92",X"06",X"6E",X"92",X"01",X"4E",X"92",X"01",X"53",X"92",X"06",X"2E",X"92",X"06",X"0E",X"92",
		X"06",X"CE",X"91",X"06",X"AE",X"91",X"02",X"8F",X"91",X"02",X"71",X"91",X"06",X"4E",X"91",X"06",
		X"0E",X"91",X"06",X"EE",X"90",X"01",X"CE",X"90",X"01",X"D1",X"90",X"01",X"D3",X"90",X"02",X"AE",
		X"90",X"03",X"B1",X"90",X"02",X"8E",X"90",X"02",X"91",X"90",X"00",X"C2",X"BC",X"48",X"3A",X"01",
		X"6B",X"A7",X"C2",X"BC",X"48",X"C3",X"97",X"49",X"C2",X"C9",X"48",X"3A",X"01",X"6B",X"A7",X"C2",
		X"C9",X"48",X"C3",X"9D",X"49",X"CD",X"F0",X"45",X"C3",X"EB",X"47",X"CD",X"C0",X"47",X"21",X"8C",
		X"38",X"C9",X"3E",X"40",X"CD",X"78",X"42",X"E1",X"23",X"23",X"3E",X"44",X"CD",X"78",X"42",X"E1",
		X"01",X"00",X"0C",X"09",X"E5",X"3E",X"17",X"CD",X"89",X"42",X"E1",X"23",X"23",X"C3",X"FC",X"45",
		X"21",X"5C",X"38",X"CD",X"32",X"3F",X"3E",X"01",X"32",X"00",X"A0",X"21",X"72",X"69",X"0E",X"6B",
		X"FF",X"21",X"73",X"69",X"0E",X"70",X"FF",X"3E",X"03",X"C3",X"20",X"52",X"21",X"CB",X"38",X"22",
		X"C4",X"63",X"3E",X"09",X"CD",X"F0",X"51",X"2A",X"C4",X"63",X"7E",X"FE",X"7F",X"CA",X"A0",X"52",
		X"23",X"22",X"C4",X"63",X"21",X"73",X"69",X"4F",X"FF",X"21",X"72",X"69",X"0E",X"FF",X"FF",X"C3",
		X"22",X"50",X"3E",X"00",X"32",X"07",X"60",X"3E",X"03",X"32",X"82",X"60",X"3E",X"F0",X"CD",X"F0",
		X"51",X"21",X"02",X"6B",X"35",X"C2",X"1C",X"50",X"3E",X"24",X"32",X"80",X"69",X"3E",X"50",X"CD",
		X"F0",X"51",X"3E",X"23",X"32",X"80",X"69",X"3E",X"50",X"CD",X"F0",X"51",X"3E",X"24",X"32",X"80",
		X"69",X"3E",X"F0",X"CD",X"F0",X"51",X"CD",X"20",X"54",X"00",X"C3",X"D4",X"53",X"FF",X"FF",X"8A",
		X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"87",X"88",X"89",X"FD",X"FD",X"FD",X"FD",X"84",X"85",X"86",
		X"FF",X"FF",X"FF",X"FF",X"81",X"82",X"83",X"FF",X"FD",X"FD",X"FF",X"80",X"FD",X"FD",X"FF",X"14",
		X"15",X"FF",X"FD",X"FD",X"FD",X"FF",X"16",X"17",X"FF",X"FD",X"FD",X"FD",X"FF",X"10",X"11",X"FF",
		X"FD",X"FD",X"FD",X"FF",X"12",X"13",X"FF",X"FD",X"FD",X"FD",X"FF",X"0C",X"0D",X"FF",X"FD",X"FD",
		X"FD",X"FF",X"0E",X"0F",X"FF",X"FD",X"FD",X"FD",X"FF",X"08",X"09",X"FF",X"FD",X"FD",X"FD",X"FF",
		X"0A",X"0B",X"FF",X"FD",X"FD",X"FD",X"FF",X"04",X"05",X"FF",X"FD",X"FD",X"FD",X"FF",X"06",X"07",
		X"FF",X"FD",X"FD",X"FD",X"FF",X"00",X"01",X"FF",X"FD",X"FD",X"FD",X"FF",X"02",X"03",X"FF",X"FD",
		X"FD",X"FD",X"FF",X"FD",X"FD",X"FF",X"FD",X"FD",X"FD",X"FF",X"FF",X"FF",X"FF",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"32",X"32",
		X"32",X"32",X"0C",X"0C",X"0C",X"32",X"32",X"32",X"32",X"0C",X"00",X"00",X"32",X"3C",X"3C",X"32",
		X"0C",X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",
		X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",
		X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",X"3C",X"3C",
		X"32",X"00",X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",
		X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",
		X"32",X"3C",X"3C",X"32",X"00",X"00",X"00",X"32",X"32",X"32",X"32",X"FD",X"FD",X"FD",X"1D",X"1E",
		X"1F",X"20",X"21",X"22",X"23",X"FD",X"1C",X"24",X"FD",X"FD",X"FD",X"FD",X"1C",X"25",X"26",X"27",
		X"28",X"29",X"2A",X"2B",X"FD",X"FD",X"FD",X"FD",X"1C",X"1B",X"FD",X"FD",X"FD",X"FD",X"1C",X"46",
		X"47",X"40",X"40",X"41",X"42",X"1B",X"FD",X"FD",X"FD",X"FD",X"1C",X"18",X"1A",X"1A",X"1A",X"1A",
		X"19",X"1B",X"FD",X"FD",X"FD",X"FD",X"1C",X"1B",X"FD",X"FD",X"FD",X"FD",X"1C",X"46",X"47",X"48",
		X"48",X"49",X"4A",X"1B",X"FD",X"FD",X"FD",X"FD",X"1C",X"2C",X"FD",X"FD",X"FD",X"FD",X"1C",X"2D",
		X"2E",X"2F",X"30",X"31",X"32",X"33",X"FD",X"FD",X"FD",X"FD",X"1C",X"34",X"35",X"36",X"37",X"FD",
		X"1C",X"FD",X"FD",X"FD",X"38",X"39",X"3A",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C3",X"70",X"54",X"C2",X"F2",X"51",X"3D",X"C2",X"F2",X"51",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"07",X"E5",X"DD",X"7E",X"00",X"77",X"23",X"DD",X"23",X"0D",X"20",X"F6",X"E1",X"19",X"10",
		X"EF",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"32",X"02",X"6B",X"AF",X"3E",X"20",X"CD",X"F0",X"51",X"00",X"00",X"00",X"00",X"AF",X"32",X"88",
		X"60",X"C3",X"1C",X"50",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"80",X"98",X"01",X"20",X"00",X"ED",X"B0",X"C9",X"FF",X"FF",X"CD",X"C0",X"53",X"C9",X"FF",
		X"0E",X"07",X"E5",X"77",X"23",X"0D",X"20",X"FB",X"E1",X"19",X"10",X"F4",X"C9",X"FF",X"FF",X"FF",
		X"11",X"20",X"00",X"21",X"49",X"9D",X"06",X"0B",X"E5",X"77",X"23",X"77",X"E1",X"19",X"10",X"F8",
		X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"C5",X"90",X"11",X"20",X"00",X"06",X"12",X"00",X"DD",X"21",X"7F",X"50",X"CD",X"00",X"52",
		X"21",X"C5",X"9C",X"DD",X"21",X"FD",X"50",X"06",X"12",X"CD",X"00",X"52",X"C9",X"FF",X"FF",X"FF",
		X"3A",X"49",X"9D",X"FE",X"3C",X"CA",X"B5",X"52",X"FE",X"31",X"CA",X"B9",X"52",X"3E",X"30",X"CD",
		X"60",X"52",X"C3",X"42",X"50",X"3E",X"31",X"18",X"F6",X"3E",X"35",X"18",X"F2",X"FF",X"FF",X"FF",
		X"21",X"C5",X"90",X"11",X"20",X"00",X"06",X"12",X"00",X"3E",X"FD",X"CD",X"50",X"52",X"21",X"C5",
		X"9C",X"3E",X"00",X"06",X"12",X"CD",X"50",X"52",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"06",X"0E",X"36",X"B0",X"23",X"10",X"FB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"20",X"00",X"06",X"0E",X"36",X"B0",X"19",X"10",X"FB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"0C",X"91",X"CD",X"E0",X"52",X"21",X"EC",X"92",X"CD",X"E0",X"52",X"21",X"2C",X"91",X"CD",
		X"F0",X"52",X"21",X"39",X"91",X"CD",X"F0",X"52",X"CD",X"20",X"53",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"21",X"0C",X"9D",X"11",X"20",X"00",X"06",X"10",X"00",X"0E",X"0E",X"E5",X"36",X"02",X"0D",X"23",
		X"20",X"FA",X"E1",X"19",X"10",X"F3",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"0C",X"91",X"11",X"20",X"00",X"06",X"10",X"0E",X"0E",X"E5",X"36",X"FD",X"23",X"0D",X"20",
		X"FA",X"E1",X"19",X"10",X"F3",X"CD",X"F0",X"45",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",
		X"21",X"FA",X"90",X"11",X"20",X"00",X"06",X"12",X"DD",X"21",X"7B",X"51",X"CD",X"00",X"5A",X"CD",
		X"80",X"53",X"C9",X"32",X"07",X"60",X"3E",X"04",X"32",X"8A",X"60",X"3D",X"32",X"1B",X"60",X"C9",
		X"21",X"FA",X"9C",X"11",X"20",X"00",X"06",X"12",X"0E",X"06",X"E5",X"36",X"34",X"23",X"0D",X"20",
		X"FA",X"E1",X"19",X"10",X"F3",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"FA",X"90",X"11",X"20",X"00",X"06",X"12",X"0E",X"06",X"E5",X"36",X"FD",X"23",X"0D",X"20",
		X"FA",X"E1",X"19",X"10",X"F3",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"30",X"54",X"CD",X"80",X"52",X"CD",X"00",
		X"53",X"C3",X"00",X"50",X"CD",X"55",X"53",X"CD",X"60",X"53",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"00",X"32",X"07",X"60",X"3E",X"04",X"32",X"8A",X"60",X"3E",X"03",X"32",X"8B",X"60",X"C3",
		X"90",X"54",X"CD",X"40",X"53",X"CD",X"A0",X"53",X"CD",X"C0",X"52",X"FD",X"E1",X"DD",X"E1",X"E1",
		X"D1",X"C1",X"F1",X"C9",X"21",X"D1",X"40",X"11",X"F3",X"4C",X"3E",X"1A",X"C3",X"51",X"54",X"FF",
		X"3E",X"00",X"32",X"07",X"60",X"3E",X"03",X"32",X"82",X"60",X"21",X"1A",X"60",X"C9",X"FF",X"FF",
		X"AF",X"32",X"07",X"60",X"3E",X"04",X"32",X"8A",X"60",X"3D",X"32",X"8B",X"60",X"C9",X"FF",X"FF",
		X"21",X"DD",X"98",X"36",X"07",X"23",X"36",X"4D",X"23",X"36",X"50",X"21",X"30",X"88",X"11",X"20",
		X"00",X"06",X"07",X"0E",X"0C",X"E5",X"36",X"A4",X"23",X"0D",X"20",X"FA",X"E1",X"19",X"10",X"F3",
		X"C9",X"A7",X"84",X"67",X"7A",X"C6",X"1F",X"57",X"7E",X"12",X"C3",X"02",X"55",X"FF",X"FF",X"FF",
		X"AF",X"0E",X"09",X"CD",X"F0",X"51",X"0D",X"C2",X"63",X"54",X"C3",X"E0",X"53",X"32",X"FF",X"6B",
		X"06",X"00",X"F5",X"3A",X"05",X"60",X"FE",X"02",X"CA",X"85",X"54",X"F1",X"05",X"C2",X"72",X"54",
		X"3D",X"C2",X"72",X"54",X"C9",X"F1",X"33",X"33",X"C3",X"FB",X"53",X"CD",X"F0",X"45",X"C9",X"FF",
		X"AF",X"0E",X"05",X"CD",X"F0",X"51",X"0D",X"C2",X"93",X"54",X"C3",X"F2",X"53",X"FF",X"FF",X"FF",
		X"10",X"10",X"10",X"FF",X"0F",X"00",X"40",X"0B",X"01",X"0B",X"01",X"0B",X"01",X"10",X"FD",X"00",
		X"FD",X"00",X"FD",X"00",X"20",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"20",X"E0",X"00",X"E0",X"00",
		X"E0",X"00",X"20",X"D5",X"00",X"D5",X"00",X"D5",X"00",X"20",X"C9",X"00",X"C9",X"00",X"C9",X"00",
		X"20",X"BD",X"00",X"BD",X"00",X"BD",X"00",X"20",X"C9",X"00",X"C9",X"00",X"C9",X"00",X"20",X"D5",
		X"00",X"D5",X"00",X"D5",X"00",X"20",X"E0",X"00",X"E0",X"00",X"E0",X"00",X"10",X"F0",X"00",X"F0",
		X"00",X"F0",X"00",X"10",X"FD",X"00",X"FD",X"00",X"FD",X"00",X"FF",X"0B",X"01",X"0B",X"01",X"0B",
		X"01",X"00",X"1B",X"23",X"23",X"7E",X"12",X"C3",X"D5",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"AF",X"32",X"FF",X"6B",
		X"CD",X"C0",X"47",X"CD",X"74",X"08",X"CD",X"C0",X"53",X"3E",X"01",X"32",X"07",X"60",X"AF",X"32",
		X"FF",X"6B",X"32",X"00",X"A0",X"32",X"0A",X"60",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"00",X"32",X"88",X"69",X"3E",X"19",X"32",X"89",X"69",X"C3",X"F8",X"18",X"3A",X"09",X"60",
		X"A7",X"C2",X"4C",X"55",X"2A",X"75",X"08",X"EB",X"2A",X"8F",X"08",X"2E",X"79",X"19",X"11",X"F2",
		X"6B",X"7E",X"12",X"6F",X"3E",X"21",X"85",X"6F",X"13",X"7E",X"12",X"C3",X"4C",X"55",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"F2",X"6B",X"A7",X"C2",X"D5",X"08",X"C3",X"04",X"54",
		X"11",X"20",X"00",X"21",X"8B",X"90",X"3E",X"FD",X"77",X"19",X"77",X"2E",X"93",X"CD",X"37",X"57",
		X"2E",X"9B",X"CD",X"37",X"57",X"21",X"4F",X"93",X"CD",X"37",X"57",X"2E",X"57",X"CD",X"37",X"57",
		X"3A",X"29",X"62",X"FE",X"01",X"28",X"0C",X"21",X"2E",X"91",X"3E",X"FD",X"77",X"21",X"12",X"92",
		X"77",X"2C",X"77",X"21",X"DC",X"3D",X"C9",X"77",X"2C",X"77",X"19",X"77",X"2D",X"77",X"C9",X"FF",
		X"3A",X"29",X"62",X"FE",X"01",X"28",X"0C",X"CB",X"7E",X"3E",X"FE",X"C2",X"F8",X"26",X"3E",X"02",
		X"C3",X"F8",X"26",X"CB",X"7E",X"3E",X"FF",X"C3",X"F3",X"26",X"CD",X"1C",X"01",X"C3",X"E7",X"57",
		X"3A",X"29",X"62",X"FE",X"01",X"28",X"11",X"21",X"D1",X"92",X"3E",X"FD",X"77",X"21",X"DD",X"91",
		X"77",X"21",X"57",X"90",X"77",X"2E",X"5A",X"77",X"21",X"00",X"62",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"2C",X"77",X"3A",X"27",X"62",X"FE",X"04",X"C0",X"3A",X"83",X"98",X"FE",X"4A",X"D0",X"3A",X"72",
		X"69",X"FE",X"62",X"D8",X"FE",X"9E",X"D0",X"AF",X"32",X"00",X"62",X"C9",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"00",X"21",X"45",X"9C",X"11",X"10",X"00",X"0E",X"1B",X"06",X"10",X"77",X"23",X"10",X"FC",
		X"19",X"0D",X"20",X"F6",X"3A",X"8A",X"63",X"C9",X"3E",X"0A",X"32",X"F7",X"9E",X"C3",X"5A",X"57",
		X"21",X"50",X"91",X"11",X"00",X"58",X"CD",X"D3",X"57",X"21",X"50",X"9D",X"CD",X"D3",X"57",X"21",
		X"88",X"63",X"C9",X"0E",X"0C",X"06",X"06",X"1A",X"77",X"23",X"13",X"10",X"FA",X"D5",X"11",X"1A",
		X"00",X"19",X"D1",X"0D",X"20",X"EF",X"C9",X"A7",X"7C",X"D6",X"1B",X"67",X"3E",X"1F",X"85",X"6F",
		X"7E",X"0F",X"0F",X"D0",X"23",X"2C",X"7E",X"0F",X"0F",X"D0",X"C3",X"F3",X"59",X"FF",X"FF",X"FF",
		X"4A",X"FD",X"FD",X"FD",X"FD",X"FD",X"FD",X"4A",X"FD",X"FD",X"FD",X"FD",X"36",X"FD",X"4A",X"4B",
		X"FD",X"FD",X"20",X"FD",X"FD",X"FD",X"4A",X"FD",X"25",X"FD",X"FD",X"FD",X"FD",X"4A",X"FD",X"FD",
		X"FD",X"FD",X"FD",X"FD",X"15",X"FD",X"FD",X"FD",X"FD",X"FD",X"26",X"FD",X"FD",X"FD",X"FD",X"48",
		X"19",X"FD",X"FD",X"FD",X"48",X"FD",X"17",X"FD",X"48",X"49",X"FD",X"FD",X"FD",X"48",X"FD",X"FD",
		X"FD",X"FD",X"48",X"FD",X"FD",X"FD",X"FD",X"FD",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"0C",X"22",X"22",X"22",X"22",X"22",X"0C",X"22",X"22",X"22",X"22",X"22",
		X"0C",X"22",X"22",X"22",X"22",X"22",X"0C",X"22",X"22",X"22",X"22",X"22",X"0C",X"22",X"22",X"22",
		X"22",X"22",X"0C",X"22",X"22",X"22",X"22",X"22",X"0C",X"22",X"22",X"22",X"22",X"22",X"0C",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"76",X"91",X"11",X"30",X"59",X"CD",X"12",X"59",X"21",X"76",X"9D",X"CD",X"12",X"59",X"C3",
		X"A0",X"57",X"0E",X"0A",X"06",X"05",X"1A",X"77",X"23",X"13",X"10",X"FA",X"D5",X"11",X"1B",X"00",
		X"19",X"D1",X"0D",X"20",X"EF",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"B0",X"B0",X"B0",X"B0",X"B0",X"B0",X"FD",X"FD",X"FD",X"B0",X"B0",X"FD",X"33",X"FD",X"B0",X"B0",
		X"FD",X"FD",X"FD",X"B0",X"B0",X"FD",X"24",X"FD",X"B0",X"B0",X"FD",X"22",X"FD",X"B0",X"B0",X"FD",
		X"11",X"FD",X"B0",X"B0",X"FD",X"20",X"FD",X"B0",X"B0",X"FD",X"FD",X"FD",X"B0",X"B0",X"B0",X"B0",
		X"B0",X"B0",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"01",X"02",
		X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"01",X"02",X"02",
		X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"02",X"02",X"01",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"03",X"92",X"11",X"1C",X"00",X"0E",X"02",X"3E",X"FD",X"06",X"04",X"77",X"23",X"10",X"FC",
		X"19",X"0D",X"20",X"F6",X"C3",X"6F",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"21",X"05",X"9D",X"06",X"03",X"77",X"23",X"10",X"FC",X"21",X"E3",X"9E",X"11",X"40",X"00",
		X"3E",X"0C",X"06",X"04",X"77",X"19",X"10",X"FC",X"C3",X"D5",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3E",X"0D",X"32",X"8A",X"60",X"01",X"E0",X"0B",X"C3",X"78",X"44",X"3E",X"0D",X"32",X"8A",X"60",
		X"C3",X"7F",X"44",X"2E",X"F2",X"3E",X"09",X"84",X"67",X"EB",X"1A",X"6F",X"13",X"1A",X"67",X"E9",
		X"0E",X"06",X"E5",X"DD",X"7E",X"00",X"77",X"23",X"DD",X"23",X"0D",X"20",X"F6",X"E1",X"19",X"10",
		X"EF",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0E",X"0B",X"E5",X"06",X"1C",X"79",X"87",X"CD",X"61",X"4A",X"5E",X"23",X"56",X"DD",X"7E",X"00",
		X"DD",X"23",X"EB",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"E1",X"0D",X"20",X"E4",X"C9",X"FF",
		X"DD",X"E5",X"21",X"6E",X"5A",X"DD",X"21",X"86",X"5A",X"CD",X"20",X"5A",X"DD",X"E1",X"21",X"8C",
		X"92",X"11",X"01",X"02",X"C9",X"FF",X"FF",X"FF",X"DD",X"E5",X"21",X"8F",X"5A",X"DD",X"21",X"A7",
		X"5A",X"CD",X"20",X"5A",X"DD",X"E1",X"C9",X"CD",X"58",X"5A",X"00",X"00",X"00",X"C3",X"B2",X"5A",
		X"47",X"9C",X"4A",X"9C",X"4C",X"9C",X"4E",X"9C",X"52",X"9C",X"54",X"9C",X"56",X"9C",X"58",X"9C",
		X"5A",X"9C",X"5C",X"9C",X"5F",X"9C",X"01",X"03",X"0B",X"02",X"0C",X"00",X"01",X"02",X"05",X"0C",
		X"00",X"47",X"9C",X"49",X"9C",X"4C",X"9C",X"4E",X"9C",X"52",X"9C",X"54",X"9C",X"56",X"9C",X"58",
		X"9C",X"5A",X"9C",X"5C",X"9C",X"5F",X"9C",X"01",X"03",X"0B",X"02",X"0C",X"00",X"01",X"02",X"05",
		X"0C",X"00",X"3A",X"0A",X"60",X"EF",X"BA",X"08",X"F8",X"08",X"21",X"1D",X"92",X"11",X"D0",X"5A",
		X"06",X"06",X"1A",X"77",X"D5",X"11",X"20",X"00",X"19",X"D1",X"13",X"10",X"F5",X"C3",X"00",X"59",
		X"1E",X"1F",X"13",X"1C",X"11",X"16",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
