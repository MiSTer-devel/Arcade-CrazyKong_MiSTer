library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_tile_bit0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_tile_bit0 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C2",X"82",X"86",X"7C",X"38",X"00",X"02",X"02",X"FE",X"FE",X"42",X"02",X"00",X"00",
		X"62",X"F2",X"BA",X"9A",X"9E",X"CE",X"46",X"00",X"8C",X"DE",X"F2",X"B2",X"92",X"86",X"04",X"00",
		X"08",X"FE",X"FE",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BE",X"A2",X"A2",X"A2",X"E6",X"E4",X"00",
		X"0C",X"9E",X"92",X"92",X"D2",X"7E",X"3C",X"00",X"C0",X"E0",X"B0",X"9E",X"8E",X"C0",X"C0",X"00",
		X"0C",X"6E",X"9A",X"9A",X"B2",X"F2",X"6C",X"00",X"78",X"FC",X"96",X"92",X"92",X"F2",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"24",X"42",X"D5",X"AB",X"42",X"24",X"18",X"00",X"00",X"80",X"80",X"80",X"80",X"FF",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"7E",X"C8",X"88",X"C8",X"7E",X"3E",X"00",
		X"6C",X"FE",X"92",X"92",X"92",X"FE",X"FE",X"00",X"44",X"C6",X"82",X"82",X"C6",X"7C",X"38",X"00",
		X"38",X"7C",X"C6",X"82",X"82",X"FE",X"FE",X"00",X"82",X"92",X"92",X"92",X"FE",X"FE",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FE",X"FE",X"00",X"9E",X"9E",X"92",X"82",X"C6",X"7C",X"38",X"00",
		X"FE",X"FE",X"10",X"10",X"10",X"FE",X"FE",X"00",X"82",X"82",X"FE",X"FE",X"82",X"82",X"00",X"00",
		X"FC",X"FE",X"02",X"02",X"02",X"06",X"04",X"00",X"82",X"C6",X"6E",X"3C",X"18",X"FE",X"FE",X"00",
		X"02",X"02",X"02",X"02",X"FE",X"FE",X"00",X"00",X"FE",X"FE",X"70",X"38",X"70",X"FE",X"FE",X"00",
		X"FE",X"FE",X"1C",X"38",X"70",X"FE",X"FE",X"00",X"7C",X"FE",X"82",X"82",X"82",X"FE",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FE",X"FE",X"00",X"7A",X"FC",X"8E",X"8A",X"82",X"FE",X"7C",X"00",
		X"72",X"F6",X"9E",X"8C",X"88",X"FE",X"FE",X"00",X"0C",X"5E",X"D2",X"92",X"92",X"F6",X"64",X"00",
		X"80",X"80",X"FE",X"FE",X"80",X"80",X"00",X"00",X"FC",X"FE",X"02",X"02",X"02",X"FE",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0E",X"1C",X"F8",X"F0",X"00",X"F8",X"FE",X"1C",X"38",X"1C",X"FE",X"F8",X"00",
		X"C6",X"EE",X"7C",X"38",X"7C",X"EE",X"C6",X"00",X"C0",X"F0",X"1E",X"1E",X"F0",X"C0",X"00",X"00",
		X"C2",X"E2",X"F2",X"BA",X"9E",X"8E",X"86",X"00",X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"00",X"00",X"28",X"00",X"00",X"00",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",
		X"00",X"00",X"82",X"C6",X"6C",X"38",X"00",X"00",X"00",X"00",X"38",X"6C",X"C6",X"82",X"00",X"00",
		X"00",X"00",X"82",X"FE",X"FE",X"82",X"00",X"00",X"82",X"FE",X"FE",X"82",X"82",X"FE",X"FE",X"82",
		X"00",X"28",X"28",X"28",X"28",X"28",X"28",X"00",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"F6",X"F6",X"00",X"00",X"F6",X"F6",X"00",X"00",X"FA",X"FA",X"00",X"00",X"FA",X"FA",X"00",X"00",
		X"00",X"00",X"00",X"F6",X"F6",X"00",X"00",X"00",X"00",X"00",X"00",X"FA",X"FA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E0",X"C0",X"00",X"00",X"00",X"00",X"E0",X"C0",X"00",X"E0",X"C0",X"00",X"00",
		X"00",X"60",X"E0",X"00",X"60",X"E0",X"00",X"00",X"00",X"00",X"C0",X"00",X"C0",X"00",X"00",X"00",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"06",X"00",X"00",
		X"38",X"28",X"3E",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"3C",X"02",X"02",X"3C",X"00",X"0E",
		X"22",X"2A",X"3E",X"00",X"00",X"0E",X"3A",X"2A",X"22",X"3E",X"00",X"3E",X"08",X"10",X"3E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"22",X"A5",X"BD",X"81",X"42",X"3C",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"42",X"81",X"A5",X"FE",X"C2",X"82",X"BA",X"44",X"44",X"28",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"0C",X"08",X"84",X"FC",X"FC",X"FC",X"FC",
		X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FB",X"F8",X"78",X"5E",X"4E",X"4E",X"40",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"03",X"07",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A3",X"59",X"FD",X"FD",X"9D",X"8C",X"88",X"00",X"00",X"00",X"01",X"03",X"31",X"59",X"28",X"5C",
		X"00",X"00",X"00",X"00",X"80",X"78",X"FC",X"7F",X"00",X"00",X"07",X"0F",X"0E",X"09",X"07",X"00",
		X"40",X"A0",X"50",X"B0",X"D0",X"68",X"B8",X"50",X"3E",X"9E",X"AE",X"DA",X"CA",X"DE",X"CD",X"D1",
		X"3F",X"7B",X"F1",X"FB",X"7F",X"FF",X"FD",X"78",X"00",X"0C",X"1E",X"3F",X"3F",X"3E",X"3E",X"1C",
		X"B8",X"50",X"A8",X"50",X"B0",X"50",X"A0",X"40",X"D1",X"D1",X"CD",X"DE",X"DA",X"AA",X"BE",X"9E",
		X"7D",X"7F",X"FF",X"FE",X"7C",X"FE",X"7F",X"3F",X"1E",X"3C",X"3E",X"3E",X"3F",X"1E",X"0C",X"00",
		X"00",X"88",X"8C",X"9D",X"FD",X"FD",X"59",X"A3",X"AE",X"1C",X"6D",X"19",X"33",X"01",X"00",X"00",
		X"7F",X"FF",X"7E",X"BE",X"1C",X"00",X"00",X"00",X"00",X"07",X"09",X"0E",X"0F",X"07",X"00",X"00",
		X"45",X"07",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"BE",X"BC",X"F8",X"E0",X"C0",X"C0",X"E0",X"03",X"01",X"01",X"03",X"07",X"0F",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"C0",X"F3",X"E2",X"C4",X"07",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"A8",X"E8",X"F9",X"FB",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"FC",X"FE",X"FF",X"FF",X"FE",X"FF",X"FE",X"AA",X"AA",X"AA",X"AA",X"EA",X"FA",X"FE",X"FF",
		X"00",X"80",X"80",X"A0",X"A0",X"A0",X"A8",X"A8",X"01",X"01",X"03",X"07",X"0F",X"1F",X"1F",X"7F",
		X"80",X"80",X"80",X"A0",X"A0",X"A8",X"A8",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"C0",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"7F",X"80",X"80",X"80",X"00",X"00",
		X"20",X"20",X"20",X"20",X"C0",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"7F",X"00",X"00",X"00",
		X"00",X"7F",X"40",X"40",X"40",X"40",X"40",X"40",X"00",X"FE",X"02",X"02",X"02",X"02",X"02",X"02",
		X"40",X"40",X"40",X"40",X"40",X"40",X"7F",X"00",X"02",X"02",X"02",X"02",X"02",X"02",X"FE",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"01",X"04",X"0E",X"8C",X"CC",X"EE",X"EE",X"EE",X"EE",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"EC",X"6C",X"0E",X"0E",X"0E",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"02",X"00",X"00",X"00",X"00",X"DE",X"3E",X"7E",X"7E",
		X"02",X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"7E",X"7E",X"7E",X"3E",X"DE",X"00",X"00",X"00",
		X"07",X"0F",X"1E",X"3F",X"3F",X"7F",X"7E",X"7E",X"80",X"00",X"00",X"00",X"80",X"00",X"04",X"02",
		X"7F",X"7E",X"7F",X"3F",X"3F",X"1E",X"0F",X"07",X"FC",X"00",X"00",X"80",X"00",X"00",X"00",X"80",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FE",
		X"1F",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"00",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",
		X"0F",X"1F",X"3F",X"3F",X"3F",X"3F",X"1D",X"08",X"00",X"C0",X"E0",X"F0",X"F0",X"F8",X"F4",X"E0",
		X"02",X"17",X"3F",X"3F",X"3F",X"3F",X"1F",X"0F",X"4A",X"1C",X"B8",X"F0",X"F0",X"E0",X"C0",X"00",
		X"00",X"01",X"0D",X"1C",X"61",X"C9",X"ED",X"C7",X"38",X"BC",X"9C",X"DC",X"FC",X"BC",X"F8",X"F8",
		X"C7",X"ED",X"C9",X"61",X"9C",X"0D",X"01",X"00",X"F8",X"FC",X"BE",X"FE",X"DE",X"8C",X"8C",X"00",
		X"03",X"07",X"05",X"08",X"1B",X"19",X"05",X"3F",X"E0",X"F0",X"50",X"08",X"6C",X"CC",X"A0",X"FE",
		X"3F",X"0F",X"05",X"37",X"3F",X"3F",X"3E",X"1C",X"FE",X"F8",X"D0",X"FB",X"FF",X"FF",X"3E",X"0C",
		X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"7E",X"42",X"42",X"42",X"42",X"42",X"42",X"7E",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"41",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"41",
		X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"FF",X"F7",X"FF",X"F7",X"F7",X"FF",X"F7",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"7F",X"80",X"F7",X"FF",X"F7",X"F7",X"FF",X"01",X"FE",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"5E",X"3F",X"07",X"05",X"09",X"7B",X"01",X"3D",
		X"06",X"0C",X"0E",X"0F",X"0F",X"07",X"03",X"00",X"7F",X"7F",X"BF",X"FF",X"FF",X"F0",X"F8",X"70",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"08",X"08",X"07",X"00",X"00",X"0F",X"04",X"00",X"20",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"FF",
		X"7F",X"44",X"44",X"44",X"44",X"44",X"44",X"7F",X"3F",X"24",X"24",X"24",X"24",X"24",X"24",X"3F",
		X"1F",X"14",X"14",X"14",X"14",X"14",X"14",X"1F",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0F",
		X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"07",X"83",X"82",X"82",X"82",X"82",X"82",X"82",X"83",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"08",X"0D",X"0B",X"09",X"08",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"20",X"00",
		X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"A0",X"20",X"20",X"20",X"20",X"20",X"20",X"A0",
		X"D0",X"50",X"50",X"50",X"50",X"50",X"50",X"D0",X"E8",X"48",X"48",X"48",X"48",X"48",X"48",X"E8",
		X"F4",X"44",X"44",X"44",X"44",X"44",X"44",X"F4",X"FA",X"42",X"42",X"42",X"42",X"42",X"42",X"FA",
		X"FD",X"45",X"45",X"45",X"45",X"45",X"45",X"FD",X"FE",X"44",X"44",X"44",X"44",X"44",X"44",X"FE",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"09",X"0A",X"0A",X"0A",X"0E",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"40",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"00",X"C0",X"00",X"C0",X"20",X"20",X"20",X"C0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"40",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"00",X"01",X"03",X"01",X"06",X"0D",X"05",X"07",X"E0",X"F0",X"F0",X"F0",X"F0",X"70",X"F0",X"F0",
		X"02",X"07",X"02",X"02",X"01",X"01",X"00",X"00",X"F0",X"70",X"F0",X"F0",X"70",X"F0",X"F0",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"F0",X"00",X"F0",X"40",X"40",X"E0",X"E0",
		X"00",X"04",X"04",X"FC",X"F8",X"00",X"A8",X"A8",X"E0",X"F8",X"7D",X"01",X"70",X"88",X"FE",X"FE",
		X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"81",X"00",X"00",X"18",X"18",X"00",X"00",X"81",X"24",X"6D",X"CF",X"EE",X"8E",X"DF",X"51",X"00",
		X"00",X"00",X"12",X"01",X"00",X"22",X"00",X"02",X"00",X"00",X"14",X"64",X"EB",X"03",X"94",X"A7",
		X"40",X"10",X"02",X"00",X"00",X"00",X"00",X"00",X"6F",X"35",X"05",X"2A",X"30",X"0C",X"02",X"00",
		X"00",X"01",X"00",X"20",X"00",X"43",X"10",X"00",X"00",X"80",X"F6",X"38",X"0F",X"3D",X"CF",X"84",
		X"00",X"40",X"21",X"02",X"00",X"00",X"00",X"00",X"5B",X"07",X"01",X"8F",X"7C",X"38",X"08",X"00",
		X"80",X"0A",X"75",X"1A",X"09",X"04",X"2F",X"50",X"0C",X"13",X"3D",X"F4",X"C9",X"07",X"1C",X"18",
		X"9C",X"0E",X"06",X"35",X"4A",X"07",X"00",X"20",X"70",X"9E",X"23",X"04",X"EC",X"9E",X"25",X"CC",
		X"08",X"80",X"00",X"00",X"09",X"86",X"40",X"01",X"00",X"0D",X"04",X"FE",X"83",X"0E",X"BC",X"BC",
		X"02",X"14",X"09",X"00",X"01",X"A6",X"43",X"00",X"78",X"9C",X"8F",X"87",X"7B",X"9D",X"01",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"7C",X"7C",X"7C",X"7C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7C",X"7C",X"7C",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"02",X"02",X"02",X"02",X"02",X"03",
		X"07",X"04",X"04",X"04",X"04",X"04",X"04",X"07",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",
		X"1F",X"11",X"11",X"11",X"11",X"11",X"11",X"1F",X"3F",X"22",X"22",X"22",X"22",X"22",X"22",X"3F",
		X"7F",X"44",X"44",X"44",X"44",X"44",X"44",X"7F",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",
		X"18",X"24",X"62",X"51",X"85",X"46",X"24",X"18",X"18",X"24",X"46",X"89",X"91",X"62",X"24",X"18",
		X"18",X"2C",X"52",X"A9",X"D5",X"4A",X"34",X"18",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"40",X"C0",X"40",X"40",X"C0",X"40",X"40",X"FF",
		X"FF",X"40",X"40",X"C0",X"40",X"40",X"C0",X"40",X"20",X"E0",X"20",X"20",X"E0",X"20",X"20",X"FF",
		X"FF",X"20",X"20",X"E0",X"20",X"20",X"E0",X"20",X"10",X"F0",X"10",X"10",X"F0",X"10",X"10",X"FF",
		X"FF",X"10",X"10",X"F0",X"10",X"10",X"F0",X"10",X"08",X"F8",X"08",X"08",X"F8",X"08",X"08",X"FF",
		X"FF",X"08",X"08",X"F8",X"08",X"08",X"F8",X"08",X"04",X"FC",X"04",X"04",X"FC",X"04",X"04",X"FF",
		X"FF",X"04",X"04",X"FC",X"04",X"04",X"FC",X"04",X"02",X"FE",X"02",X"02",X"FE",X"02",X"02",X"FF",
		X"FF",X"02",X"02",X"FE",X"02",X"02",X"FE",X"02",X"81",X"FF",X"81",X"81",X"FF",X"81",X"81",X"FF",
		X"FF",X"81",X"81",X"FF",X"81",X"81",X"FF",X"81",X"40",X"7F",X"40",X"40",X"7F",X"40",X"40",X"FF",
		X"FF",X"40",X"40",X"7F",X"40",X"40",X"7F",X"40",X"20",X"3F",X"20",X"20",X"3F",X"20",X"20",X"FF",
		X"FF",X"20",X"20",X"3F",X"20",X"20",X"3F",X"20",X"10",X"1F",X"10",X"10",X"1F",X"10",X"10",X"FF",
		X"FF",X"10",X"10",X"1F",X"10",X"10",X"1F",X"10",X"08",X"0F",X"08",X"08",X"0F",X"08",X"08",X"FF",
		X"FF",X"08",X"08",X"0F",X"08",X"08",X"0F",X"08",X"04",X"07",X"04",X"04",X"07",X"04",X"04",X"FF",
		X"FF",X"04",X"04",X"07",X"04",X"04",X"07",X"04",X"02",X"03",X"02",X"02",X"03",X"02",X"02",X"FF",
		X"FF",X"02",X"02",X"03",X"02",X"02",X"03",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"FF",
		X"FF",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"08",X"84",X"FC",X"FC",X"FC",X"FC",
		X"FB",X"F8",X"78",X"5E",X"4E",X"4E",X"40",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"07",X"0E",X"1C",X"38",X"70",X"E0",X"C0",X"83",X"87",X"8E",X"9C",X"B8",X"F0",X"E0",X"C0",
		X"C0",X"E0",X"70",X"38",X"1C",X"0E",X"07",X"03",X"C0",X"E0",X"F0",X"B8",X"9C",X"8E",X"87",X"83",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"58",X"7B",X"7F",X"1F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"67",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"A8",X"B8",X"B0",X"38",X"60",
		X"FF",X"9E",X"1C",X"0D",X"09",X"03",X"06",X"04",X"40",X"C0",X"80",X"D0",X"F0",X"E0",X"40",X"00",
		X"01",X"01",X"21",X"6C",X"FE",X"FE",X"FE",X"FF",X"80",X"40",X"E0",X"F0",X"E0",X"C0",X"40",X"40",
		X"FF",X"BF",X"DE",X"66",X"20",X"00",X"00",X"00",X"40",X"68",X"78",X"F8",X"D0",X"40",X"00",X"00",
		X"00",X"00",X"27",X"77",X"DF",X"BF",X"FF",X"FF",X"00",X"40",X"40",X"68",X"38",X"20",X"B8",X"A0",
		X"FF",X"FF",X"FF",X"5F",X"77",X"27",X"00",X"00",X"A0",X"B8",X"B0",X"38",X"68",X"40",X"40",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"44",X"44",X"44",X"44",X"44",X"44",X"FF",X"FF",X"C4",X"C4",X"C4",X"C4",X"C4",X"C4",X"FF",
		X"7F",X"44",X"44",X"44",X"44",X"44",X"44",X"7F",X"3F",X"24",X"24",X"24",X"24",X"24",X"24",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"3F",X"3F",X"00",X"00",X"00",X"E3",X"F3",X"FB",X"B9",X"10",
		X"3F",X"3F",X"1E",X"1E",X"1C",X"08",X"00",X"00",X"43",X"83",X"83",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"1D",X"3D",X"3F",X"3E",X"3E",X"E0",X"E6",X"C7",X"87",X"C1",X"C0",X"00",X"40",
		X"3F",X"3F",X"1E",X"1E",X"1C",X"09",X"01",X"00",X"00",X"80",X"80",X"C0",X"DC",X"FC",X"C0",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"1E",X"1F",X"1F",X"1E",X"1C",X"20",X"60",X"C0",X"C0",X"E0",X"E3",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0E",X"04",X"00",X"E3",X"63",X"61",X"E0",X"40",X"00",X"00",X"00",
		X"00",X"03",X"07",X"07",X"1F",X"3C",X"1F",X"1F",X"00",X"00",X"00",X"00",X"02",X"07",X"07",X"87",
		X"1F",X"1F",X"3C",X"FF",X"FF",X"1C",X"00",X"00",X"83",X"0B",X"08",X"08",X"08",X"00",X"00",X"00",
		X"00",X"10",X"30",X"20",X"40",X"60",X"70",X"70",X"00",X"00",X"00",X"00",X"06",X"0F",X"0F",X"0F",
		X"60",X"40",X"70",X"30",X"18",X"1C",X"0C",X"00",X"37",X"33",X"30",X"20",X"00",X"00",X"00",X"00",
		X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"10",X"C0",X"C0",X"00",X"00",X"0C",X"0E",X"0E",X"06",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"40",X"40",X"40",X"40",X"40",X"40",X"00",
		X"00",X"00",X"01",X"03",X"1B",X"3C",X"1F",X"1F",X"60",X"E0",X"E0",X"81",X"01",X"01",X"81",X"C1",
		X"1F",X"1F",X"3C",X"1B",X"03",X"01",X"00",X"00",X"C1",X"81",X"01",X"01",X"81",X"E0",X"E0",X"60",
		X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",X"00",X"00",X"00",X"FF",X"44",X"44",X"44",X"44",
		X"44",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",X"44",X"44",X"44",X"44",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"FF",X"FF",X"00",X"00",X"00",X"03",X"C3",X"C3",X"C1",X"80",
		X"FF",X"3E",X"1E",X"1E",X"1C",X"08",X"00",X"00",X"43",X"03",X"83",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"3F",X"3E",X"00",X"00",X"00",X"C3",X"E3",X"E3",X"C1",X"C0",
		X"3E",X"3F",X"1E",X"1E",X"1C",X"08",X"00",X"00",X"C3",X"C3",X"C3",X"C1",X"E0",X"E0",X"E0",X"C0",
		X"00",X"00",X"04",X"1C",X"3D",X"3F",X"FF",X"FF",X"00",X"06",X"07",X"03",X"C1",X"C0",X"C0",X"00",
		X"FF",X"3E",X"1E",X"1E",X"1C",X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"1C",X"3C",X"00",X"00",
		X"00",X"00",X"04",X"1C",X"3C",X"3F",X"3F",X"3E",X"00",X"06",X"07",X"03",X"C1",X"E0",X"E0",X"C0",
		X"3E",X"3F",X"1E",X"1E",X"1C",X"08",X"00",X"00",X"C0",X"C0",X"C0",X"C0",X"FC",X"FC",X"E0",X"C0",
		X"00",X"00",X"00",X"02",X"0E",X"1E",X"1F",X"FF",X"1E",X"1C",X"00",X"00",X"C0",X"C0",X"E0",X"E3",
		X"FF",X"FF",X"1F",X"0F",X"0F",X"0E",X"04",X"00",X"C3",X"A3",X"81",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"02",X"0E",X"1E",X"1F",X"1F",X"1E",X"1C",X"00",X"00",X"C0",X"C0",X"E0",X"E3",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0E",X"04",X"00",X"E3",X"63",X"E1",X"60",X"60",X"E0",X"E0",X"C0",
		X"00",X"01",X"01",X"02",X"0E",X"1E",X"1F",X"1F",X"84",X"8C",X"D8",X"9C",X"C8",X"E0",X"E0",X"00",
		X"1F",X"1F",X"1F",X"0F",X"0F",X"0E",X"05",X"01",X"20",X"80",X"C0",X"40",X"40",X"C0",X"CC",X"9C",
		X"01",X"03",X"07",X"1F",X"3F",X"3F",X"3E",X"3F",X"C1",X"E5",X"42",X"82",X"C1",X"C0",X"80",X"41",
		X"3F",X"3F",X"1F",X"1F",X"1D",X"09",X"00",X"00",X"03",X"87",X"8E",X"8D",X"83",X"C6",X"CC",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"70",X"58",X"7B",X"7F",X"1F",X"2F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"67",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"08",X"A8",X"B8",X"B0",X"38",X"60",
		X"FF",X"9E",X"1C",X"0D",X"09",X"03",X"06",X"04",X"40",X"C0",X"80",X"D0",X"F0",X"E0",X"40",X"00",
		X"01",X"01",X"21",X"6C",X"FE",X"FE",X"FE",X"FF",X"80",X"40",X"E0",X"F0",X"E0",X"C0",X"40",X"40",
		X"FF",X"BF",X"DE",X"66",X"20",X"00",X"00",X"00",X"40",X"68",X"78",X"F8",X"D0",X"40",X"00",X"00",
		X"00",X"00",X"27",X"77",X"DF",X"BF",X"FF",X"FF",X"00",X"40",X"40",X"68",X"38",X"20",X"B8",X"A0",
		X"FF",X"FF",X"FF",X"5F",X"77",X"27",X"00",X"00",X"A0",X"B8",X"B0",X"38",X"68",X"40",X"40",X"00",
		X"00",X"00",X"06",X"0E",X"1D",X"1B",X"1B",X"1B",X"40",X"C0",X"DC",X"FF",X"FF",X"C7",X"02",X"00",
		X"1A",X"1A",X"1B",X"0A",X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"60",X"00",
		X"00",X"00",X"03",X"04",X"08",X"0A",X"11",X"10",X"00",X"00",X"C0",X"20",X"10",X"10",X"08",X"88",
		X"10",X"16",X"0E",X"08",X"04",X"03",X"00",X"00",X"48",X"08",X"10",X"10",X"20",X"C0",X"00",X"00",
		X"02",X"0F",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"40",X"F0",X"20",X"20",X"30",X"30",X"30",X"30",
		X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"0F",X"02",X"30",X"30",X"30",X"30",X"20",X"20",X"F0",X"40",
		X"05",X"0F",X"0B",X"1B",X"13",X"13",X"13",X"13",X"A0",X"F0",X"D0",X"D8",X"C8",X"C8",X"C8",X"C8",
		X"13",X"13",X"13",X"13",X"1B",X"0B",X"0F",X"05",X"C8",X"C8",X"C8",X"C8",X"D8",X"D0",X"F0",X"A0",
		X"00",X"00",X"00",X"00",X"4F",X"7F",X"C0",X"40",X"00",X"00",X"00",X"00",X"F2",X"FE",X"03",X"02",
		X"40",X"C0",X"7F",X"4F",X"00",X"00",X"00",X"00",X"02",X"03",X"FF",X"F2",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"03",X"07",X"07",X"0F",X"0F",X"00",X"00",X"00",X"C0",X"E0",X"E0",X"F0",X"F0",
		X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"F0",X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",
		X"05",X"0F",X"0B",X"1B",X"13",X"13",X"13",X"13",X"A0",X"F0",X"D0",X"D8",X"C8",X"C8",X"C8",X"C8",
		X"13",X"13",X"13",X"13",X"1B",X"0B",X"0F",X"05",X"C8",X"C8",X"C8",X"C8",X"D8",X"D0",X"F0",X"A0",
		X"02",X"0F",X"04",X"04",X"0C",X"0C",X"0C",X"0C",X"40",X"F0",X"20",X"20",X"30",X"30",X"30",X"30",
		X"0C",X"0C",X"0C",X"0C",X"04",X"04",X"0F",X"02",X"30",X"30",X"30",X"30",X"20",X"20",X"F0",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"F0",X"F0",
		X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"00",X"02",X"08",X"04",X"02",X"F8",X"FC",X"FC",
		X"03",X"03",X"03",X"01",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FA",X"02",X"0A",X"14",X"02",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"BF",X"9E",X"C1",X"33",X"39",X"78",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"E1",X"C6",X"8F",X"CF",X"E6",X"73",X"1F",X"00",X"7E",X"7E",X"7E",X"7E",X"7C",X"3D",X"19",X"03",
		X"00",X"1E",X"36",X"60",X"C0",X"CC",X"ED",X"F1",X"1F",X"27",X"47",X"43",X"43",X"43",X"43",X"43",
		X"ED",X"CC",X"C0",X"60",X"36",X"1E",X"0E",X"00",X"43",X"43",X"43",X"43",X"47",X"27",X"1F",X"1F",
		X"00",X"1E",X"36",X"60",X"C0",X"CC",X"ED",X"F1",X"6F",X"F7",X"F7",X"73",X"7B",X"7B",X"7B",X"73",
		X"ED",X"CC",X"C0",X"60",X"36",X"1E",X"0E",X"00",X"7B",X"7B",X"7B",X"73",X"F7",X"F7",X"67",X"0F",
		X"FE",X"47",X"87",X"14",X"85",X"04",X"89",X"F0",X"00",X"00",X"C0",X"C0",X"40",X"C0",X"C0",X"40",
		X"F0",X"89",X"04",X"85",X"14",X"87",X"47",X"FE",X"C0",X"40",X"C0",X"40",X"C0",X"C0",X"00",X"00",
		X"00",X"01",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"E0",X"E0",X"E0",X"E0",X"F0",X"F8",X"F8",X"F8",
		X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",X"F8",X"F4",X"F0",X"F0",X"28",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"87",X"FF",X"00",X"01",X"02",X"E4",X"F8",X"FA",X"FC",X"FC",
		X"FF",X"FF",X"FF",X"FF",X"01",X"00",X"00",X"00",X"FC",X"F8",X"FA",X"FC",X"F8",X"F8",X"30",X"20",
		X"01",X"0F",X"07",X"0F",X"07",X"23",X"13",X"09",X"C0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",
		X"51",X"31",X"11",X"01",X"01",X"03",X"01",X"01",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"00",X"11",X"1F",X"1F",X"00",X"05",X"02",X"07",X"0F",X"FF",X"FF",X"FF",
		X"1F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"00",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"F8",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"3F",X"7F",X"FF",
		X"01",X"03",X"07",X"07",X"07",X"03",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",
		X"00",X"00",X"00",X"00",X"C0",X"F8",X"FE",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"EE",X"FF",X"FC",X"F0",X"00",X"C0",X"C0",X"60",X"B0",X"40",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"78",X"00",X"CC",
		X"00",X"00",X"01",X"01",X"0F",X"1F",X"3F",X"7F",X"F8",X"FE",X"FD",X"FC",X"F9",X"F8",X"F8",X"F8",
		X"F4",X"F9",X"FD",X"FE",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"FC",X"FC",X"32",X"84",X"C3",X"F0",
		X"3F",X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"F8",X"F0",X"F0",X"A0",X"04",X"02",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"F8",X"F8",X"F0",X"E0",X"E0",X"E0",X"E0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E6",X"E2",X"E0",X"E0",X"E0",X"E6",X"FC",X"78",X"F8",X"FC",
		X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",X"00",X"01",X"07",X"3F",X"FF",X"FF",X"FF",X"FF",
		X"07",X"0F",X"0F",X"0F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3C",X"78",X"78",X"FC",X"F7",X"E3",X"E1",X"C0",X"FF",X"FF",X"3F",X"9F",X"CF",X"E3",X"C1",X"80",
		X"CC",X"4C",X"00",X"04",X"04",X"00",X"00",X"00",X"08",X"10",X"20",X"20",X"20",X"20",X"20",X"00",
		X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"60",X"F0",X"F8",X"FC",X"FC",X"FE",X"FC",X"EC",
		X"07",X"07",X"0F",X"0F",X"0F",X"0F",X"0C",X"08",X"CE",X"CE",X"C0",X"C0",X"E0",X"E0",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"0F",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"00",X"00",X"00",X"00",X"00",X"0B",X"FF",X"FF",
		X"07",X"0F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"20",X"5C",X"7F",X"FF",X"7F",X"7F",X"1F",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"FF",
		X"0F",X"07",X"01",X"00",X"00",X"00",X"00",X"00",X"FE",X"FC",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"03",X"03",X"07",X"07",X"07",X"0F",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"0F",X"07",X"07",X"0B",X"00",X"00",X"00",X"00",X"FF",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"18",X"30",X"F6",X"F7",X"F7",X"F3",X"FB",
		X"FF",X"FF",X"FF",X"7F",X"1F",X"0E",X"00",X"00",X"F9",X"FC",X"E4",X"C2",X"00",X"00",X"00",X"00",
		X"00",X"1C",X"3E",X"7F",X"FF",X"FF",X"FF",X"FE",X"00",X"00",X"00",X"00",X"90",X"30",X"70",X"F0",
		X"FE",X"FE",X"FF",X"FF",X"FE",X"FE",X"FE",X"FE",X"F0",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"08",X"04",X"00",X"00",X"00",X"00",X"80",X"49",X"2A",X"08",X"7E",X"08",X"2A",X"49",
		X"00",X"00",X"00",X"00",X"00",X"01",X"02",X"00",X"80",X"00",X"02",X"09",X"80",X"08",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"40",X"61",X"63",X"66",X"6C",X"7A",X"00",X"00",X"81",X"C3",X"E3",X"33",X"1B",X"AF",
		X"7A",X"6C",X"66",X"63",X"61",X"40",X"00",X"00",X"AF",X"1B",X"33",X"E3",X"C3",X"81",X"00",X"00",
		X"00",X"00",X"04",X"06",X"06",X"06",X"06",X"07",X"20",X"70",X"71",X"53",X"DB",X"8B",X"8B",X"FF",
		X"07",X"06",X"06",X"06",X"06",X"04",X"00",X"00",X"FF",X"8B",X"8B",X"DB",X"53",X"71",X"70",X"20",
		X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"78",X"FC",X"CC",
		X"00",X"21",X"00",X"00",X"04",X"00",X"00",X"00",X"FC",X"FC",X"CC",X"78",X"00",X"00",X"00",X"00",
		X"08",X"00",X"00",X"00",X"00",X"01",X"23",X"03",X"00",X"00",X"00",X"00",X"78",X"FC",X"FE",X"CE",
		X"05",X"01",X"02",X"00",X"10",X"02",X"00",X"00",X"FE",X"FE",X"CC",X"FC",X"78",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"30",X"30",X"30",X"00",X"00",X"00",X"00",X"C0",X"C0",X"C0",X"C0",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"C0",X"C0",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"30",X"30",X"00",X"00",X"00",X"00",X"FC",X"FC",X"C0",X"C0",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"C0",X"C0",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0C",X"0C",X"0C",
		X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"0C",X"0C",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"3C",X"30",X"30",X"00",X"00",X"00",X"00",X"3C",X"3C",X"0C",X"0C",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"0C",X"0C",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"30",X"30",X"00",X"00",X"00",X"00",X"FC",X"FC",X"0C",X"0C",
		X"30",X"30",X"3F",X"3F",X"00",X"00",X"00",X"00",X"0C",X"0C",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"30",X"C0",
		X"03",X"0C",X"3F",X"3F",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"00",X"00",X"00",X"00",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FC",
		X"00",X"00",X"01",X"0F",X"7E",X"F0",X"80",X"00",X"0F",X"3F",X"FB",X"C3",X"03",X"03",X"03",X"03",
		X"00",X"00",X"00",X"00",X"00",X"03",X"1F",X"FC",X"00",X"00",X"01",X"0F",X"7E",X"F0",X"80",X"00",
		X"07",X"3F",X"F8",X"C0",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C3",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"3F",X"FF",X"C0",X"00",
		X"00",X"00",X"03",X"FF",X"FC",X"00",X"00",X"00",X"00",X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",
		X"3F",X"FF",X"C3",X"03",X"03",X"03",X"03",X"03",X"FC",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"FC",X"FF",X"C3",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"F0",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"FF",X"3F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FC",X"FF",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"0F",X"00",
		X"03",X"03",X"03",X"03",X"03",X"C3",X"FF",X"3F",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"C0",X"E0",
		X"FC",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"7E",X"0F",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"C0",X"F8",X"3F",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",
		X"FC",X"1F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"F0",X"7E",X"0F",X"01",X"00",X"00",
		X"03",X"03",X"03",X"03",X"C3",X"FD",X"3F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"03",X"03",X"03",X"03",X"03",X"03",X"FF",X"FF",
		X"C0",X"C0",X"FF",X"FF",X"C0",X"C0",X"C0",X"C0",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"03",X"03",X"03",X"03",X"FF",X"FF",X"03",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
