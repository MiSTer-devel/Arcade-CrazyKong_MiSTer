library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ckong_samples is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ckong_samples is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"99",X"99",X"99",X"87",X"55",X"68",X"99",X"AB",X"BB",X"BA",X"85",X"33",X"68",X"99",X"9B",X"BB",
		X"BA",X"74",X"23",X"79",X"99",X"9B",X"CC",X"BB",X"94",X"12",X"59",X"A9",X"9A",X"BC",X"CB",X"94",
		X"12",X"69",X"99",X"89",X"BC",X"CC",X"B6",X"20",X"27",X"9A",X"99",X"BC",X"CD",X"B5",X"10",X"37",
		X"BA",X"98",X"9C",X"ED",X"DA",X"30",X"04",X"9B",X"A8",X"9B",X"DE",X"DA",X"50",X"03",X"8B",X"B9",
		X"79",X"DF",X"FD",X"60",X"00",X"6B",X"C9",X"77",X"BF",X"FF",X"A6",X"00",X"19",X"CB",X"86",X"9D",
		X"FF",X"D5",X"00",X"06",X"CC",X"96",X"7B",X"FF",X"FB",X"10",X"03",X"AC",X"B7",X"59",X"EF",X"FB",
		X"60",X"01",X"9C",X"C8",X"68",X"EF",X"FC",X"50",X"01",X"9E",X"C8",X"58",X"DF",X"FD",X"30",X"02",
		X"9D",X"A5",X"49",X"FF",X"FB",X"40",X"04",X"CC",X"62",X"6F",X"FF",X"F4",X"00",X"2C",X"C5",X"05",
		X"EF",X"FF",X"C0",X"04",X"D9",X"00",X"BF",X"FF",X"F0",X"01",X"DB",X"00",X"DF",X"FF",X"F0",X"01",
		X"F9",X"00",X"FF",X"CF",X"F0",X"0F",X"F0",X"0C",X"F6",X"EF",X"B0",X"0F",X"71",X"1F",X"8D",X"FF",
		X"00",X"F4",X"06",X"F5",X"EF",X"F0",X"2F",X"10",X"9B",X"7F",X"F0",X"0F",X"F0",X"0F",X"6F",X"F6",
		X"0D",X"F0",X"0F",X"7F",X"F0",X"0F",X"C0",X"5F",X"9F",X"F0",X"0F",X"00",X"FC",X"FF",X"00",X"F9",
		X"06",X"FF",X"F0",X"0F",X"60",X"BF",X"FF",X"00",X"FC",X"07",X"FF",X"F0",X"0F",X"B0",X"6F",X"FF",
		X"00",X"F1",X"0A",X"FF",X"F0",X"6F",X"00",X"FF",X"F6",X"0B",X"F0",X"0C",X"FF",X"60",X"8F",X"00",
		X"CF",X"F7",X"01",X"F0",X"0F",X"FF",X"60",X"0F",X"00",X"FF",X"F7",X"00",X"71",X"0F",X"FF",X"81",
		X"03",X"43",X"FF",X"FF",X"00",X"05",X"7F",X"FF",X"F0",X"00",X"39",X"EF",X"FF",X"93",X"01",X"69",
		X"BC",X"FD",X"D9",X"87",X"98",X"6B",X"BB",X"9A",X"9B",X"88",X"87",X"46",X"78",X"76",X"89",X"96",
		X"88",X"86",X"78",X"87",X"67",X"A6",X"79",X"69",X"99",X"89",X"99",X"88",X"98",X"9B",X"A7",X"77",
		X"8A",X"9A",X"98",X"86",X"66",X"87",X"8C",X"98",X"56",X"87",X"77",X"99",X"68",X"89",X"79",X"9A",
		X"96",X"89",X"88",X"A9",X"97",X"79",X"A9",X"88",X"A9",X"78",X"57",X"AA",X"8B",X"74",X"89",X"77",
		X"7A",X"77",X"76",X"86",X"97",X"68",X"99",X"99",X"87",X"8B",X"84",X"7A",X"98",X"A9",X"89",X"87",
		X"98",X"9A",X"7B",X"96",X"58",X"B8",X"6C",X"7B",X"68",X"8B",X"8A",X"7A",X"9B",X"75",X"97",X"B8",
		X"89",X"96",X"86",X"9A",X"98",X"79",X"96",X"97",X"A6",X"77",X"97",X"A7",X"78",X"77",X"9A",X"97",
		X"B6",X"4B",X"A9",X"87",X"96",X"87",X"79",X"AA",X"75",X"65",X"89",X"87",X"88",X"79",X"79",X"78",
		X"99",X"C9",X"98",X"BB",X"88",X"66",X"78",X"75",X"74",X"88",X"77",X"58",X"ED",X"AB",X"8B",X"98",
		X"64",X"87",X"A8",X"74",X"95",X"78",X"43",X"23",X"9C",X"FF",X"EF",X"B1",X"00",X"00",X"BF",X"FF",
		X"FF",X"B0",X"00",X"00",X"0B",X"FF",X"FF",X"FA",X"00",X"11",X"21",X"4F",X"FF",X"FB",X"C9",X"01",
		X"82",X"77",X"0F",X"FD",X"F7",X"6B",X"20",X"B4",X"2E",X"62",X"FD",X"8D",X"99",X"D0",X"0C",X"05",
		X"C2",X"96",X"8C",X"99",X"65",X"E0",X"07",X"0F",X"03",X"B0",X"D7",X"76",X"4B",X"C0",X"54",X"0F",
		X"0F",X"87",X"E6",X"C5",X"98",X"CD",X"06",X"04",X"63",X"E1",X"F3",X"F6",X"B7",X"8A",X"9F",X"FE",
		X"6F",X"0F",X"0D",X"3C",X"59",X"7B",X"69",X"A6",X"C8",X"88",X"89",X"79",X"68",X"88",X"8A",X"8A",
		X"8A",X"69",X"69",X"89",X"89",X"89",X"79",X"79",X"79",X"8A",X"7A",X"59",X"69",X"78",X"70",X"70",
		X"88",X"88",X"88",X"88",X"88",X"88",X"75",X"A8",X"B8",X"88",X"88",X"78",X"77",X"98",X"97",X"87",
		X"8C",X"0B",X"3C",X"87",X"B7",X"B7",X"67",X"9B",X"88",X"88",X"97",X"99",X"BB",X"B7",X"00",X"68",
		X"62",X"4A",X"DF",X"FF",X"FF",X"00",X"1D",X"60",X"2B",X"C2",X"4C",X"DD",X"FF",X"FF",X"00",X"5E",
		X"00",X"9C",X"40",X"B9",X"9E",X"FF",X"FF",X"00",X"78",X"05",X"B3",X"39",X"73",X"BB",X"FF",X"FF",
		X"30",X"D8",X"03",X"C5",X"0D",X"45",X"8C",X"FF",X"FF",X"F0",X"0A",X"00",X"D4",X"36",X"92",X"99",
		X"FF",X"FF",X"FF",X"0F",X"10",X"0F",X"07",X"76",X"59",X"CF",X"FF",X"FF",X"40",X"F0",X"06",X"B0",
		X"75",X"39",X"9F",X"FF",X"FF",X"F0",X"F2",X"00",X"F0",X"85",X"66",X"C9",X"FF",X"FF",X"F0",X"09",
		X"00",X"D3",X"26",X"66",X"B8",X"FF",X"FF",X"F0",X"0A",X"00",X"B6",X"18",X"56",X"C9",X"FF",X"FF",
		X"F0",X"67",X"00",X"A5",X"29",X"47",X"CA",X"FF",X"FF",X"F0",X"B4",X"00",X"96",X"1A",X"48",X"BD",
		X"FF",X"FF",X"60",X"F0",X"00",X"B4",X"08",X"7A",X"BF",X"FF",X"FF",X"00",X"F0",X"00",X"A6",X"27",
		X"CD",X"CF",X"FF",X"FF",X"00",X"50",X"00",X"68",X"A9",X"99",X"9A",X"BD",X"EF",X"BA",X"41",X"00",
		X"24",X"66",X"79",X"CD",X"EF",X"FC",X"B9",X"10",X"00",X"25",X"78",X"8B",X"EF",X"FF",X"FC",X"B4",
		X"00",X"00",X"34",X"8A",X"AD",X"FF",X"FF",X"BB",X"60",X"00",X"00",X"45",X"9C",X"CE",X"FF",X"FD",
		X"A6",X"00",X"00",X"03",X"67",X"AE",X"FF",X"FF",X"FB",X"91",X"00",X"00",X"24",X"89",X"CF",X"FF",
		X"FF",X"CB",X"40",X"00",X"01",X"47",X"9C",X"FF",X"FF",X"FC",X"B5",X"00",X"00",X"03",X"69",X"BE",
		X"FF",X"FF",X"EC",X"71",X"00",X"00",X"25",X"8B",X"DF",X"FF",X"FF",X"CB",X"20",X"00",X"02",X"47",
		X"AD",X"FF",X"FF",X"FC",X"B4",X"00",X"00",X"14",X"69",X"CE",X"FF",X"FF",X"FC",X"71",X"00",X"01",
		X"25",X"7B",X"DE",X"FF",X"FF",X"CA",X"31",X"00",X"12",X"47",X"9C",X"DF",X"FF",X"FE",X"B7",X"11",
		X"00",X"23",X"57",X"AC",X"DF",X"FF",X"FC",X"94",X"11",X"02",X"35",X"68",X"BC",X"EE",X"EF",X"EB",
		X"72",X"10",X"13",X"36",X"7A",X"BC",X"EE",X"FF",X"CA",X"62",X"10",X"23",X"57",X"9B",X"CE",X"EE",
		X"ED",X"B9",X"42",X"11",X"23",X"68",X"AB",X"DE",X"DD",X"CC",X"99",X"42",X"11",X"24",X"69",X"BC",
		X"DD",X"CC",X"BB",X"98",X"64",X"23",X"35",X"69",X"BC",X"CB",X"AA",X"99",X"88",X"87",X"65",X"56",
		X"78",X"99",X"A9",X"99",X"99",X"9A",X"BA",X"96",X"54",X"45",X"67",X"89",X"99",X"AA",X"AA",X"BB",
		X"A8",X"75",X"43",X"45",X"79",X"9A",X"AA",X"64",X"3F",X"FF",X"00",X"0F",X"F0",X"06",X"F8",X"1B",
		X"FF",X"FF",X"F0",X"09",X"B0",X"0C",X"90",X"0D",X"B9",X"FF",X"FF",X"00",X"F6",X"00",X"F3",X"08",
		X"E4",X"AF",X"FF",X"FF",X"00",X"F1",X"00",X"F0",X"0F",X"17",X"9B",X"FF",X"FF",X"00",X"F1",X"03",
		X"C0",X"4F",X"09",X"AA",X"FF",X"FF",X"00",X"F2",X"0B",X"90",X"6F",X"0B",X"97",X"FF",X"FF",X"81",
		X"F1",X"05",X"A0",X"3F",X"09",X"97",X"FF",X"FF",X"F0",X"F4",X"00",X"F1",X"0F",X"08",X"B7",X"FF",
		X"FF",X"F0",X"F8",X"01",X"F1",X"0F",X"04",X"D7",X"FF",X"FF",X"F0",X"DA",X"00",X"E4",X"0F",X"01",
		X"D6",X"FF",X"FF",X"F0",X"4A",X"00",X"F7",X"0F",X"60",X"C7",X"BF",X"FF",X"F0",X"08",X"20",X"EB",
		X"0B",X"B0",X"9A",X"8F",X"FF",X"F6",X"09",X"C0",X"5D",X"04",X"D4",X"1A",X"BD",X"FF",X"FF",X"06",
		X"E0",X"0A",X"C0",X"7F",X"04",X"EA",X"FF",X"FF",X"00",X"6B",X"00",X"F4",X"0A",X"82",X"7D",X"FF",
		X"FF",X"F0",X"0E",X"10",X"2F",X"81",X"88",X"69",X"CF",X"FF",X"F5",X"00",X"66",X"56",X"37",X"98",
		X"76",X"77",X"DF",X"FF",X"E8",X"10",X"05",X"99",X"A9",X"75",X"69",X"CC",X"CD",X"EE",X"B6",X"00",
		X"03",X"AC",X"C9",X"64",X"7B",X"DE",X"EC",X"DF",X"A3",X"00",X"16",X"AC",X"C8",X"55",X"7B",X"DC",
		X"BE",X"FE",X"30",X"05",X"BA",X"43",X"6C",X"93",X"7E",X"FF",X"FF",X"F0",X"06",X"E5",X"00",X"8F",
		X"60",X"4D",X"CC",X"FF",X"F0",X"00",X"F8",X"00",X"FA",X"06",X"B6",X"8E",X"FF",X"FF",X"00",X"89",
		X"00",X"8F",X"40",X"C9",X"1A",X"FF",X"FF",X"F0",X"0F",X"A0",X"0F",X"B0",X"5F",X"40",X"CE",X"CF",
		X"FF",X"00",X"E9",X"00",X"F9",X"07",X"F5",X"0B",X"FC",X"FF",X"F6",X"04",X"C0",X"08",X"D3",X"1D",
		X"B0",X"6F",X"EE",X"FF",X"F0",X"0F",X"C0",X"0F",X"A0",X"6F",X"40",X"CF",X"CF",X"FF",X"81",X"2E",
		X"40",X"4F",X"60",X"AF",X"20",X"EF",X"CF",X"FF",X"00",X"7D",X"00",X"9E",X"30",X"CF",X"00",X"EF",
		X"AF",X"FF",X"20",X"7D",X"00",X"6D",X"71",X"8F",X"60",X"9F",X"CE",X"FF",X"81",X"2D",X"81",X"1E",
		X"D0",X"3F",X"C0",X"4E",X"DC",X"FF",X"F0",X"09",X"F0",X"0B",X"F5",X"0A",X"F8",X"07",X"ED",X"DF",
		X"FE",X"00",X"AE",X"10",X"9F",X"61",X"9F",X"90",X"5D",X"CB",X"FF",X"F0",X"08",X"D1",X"07",X"F7",
		X"18",X"FB",X"13",X"BC",X"9C",X"FF",X"81",X"4C",X"91",X"2B",X"D6",X"4C",X"F7",X"36",X"B9",X"58",
		X"CC",X"BC",X"C8",X"34",X"89",X"64",X"9B",X"75",X"8B",X"A7",X"79",X"97",X"67",X"98",X"78",X"9A",
		X"9A",X"C9",X"54",X"79",X"75",X"6A",X"96",X"79",X"A8",X"79",X"A9",X"78",X"89",X"98",X"88",X"88",
		X"99",X"87",X"88",X"88",X"99",X"87",X"79",X"99",X"87",X"89",X"98",X"87",X"88",X"88",X"70",X"70",
		X"89",X"98",X"77",X"79",X"99",X"87",X"78",X"A9",X"87",X"78",X"A9",X"87",X"79",X"A9",X"77",X"79",
		X"B8",X"77",X"79",X"A9",X"77",X"77",X"9A",X"87",X"77",X"79",X"B9",X"66",X"88",X"9B",X"B8",X"55",
		X"78",X"99",X"BB",X"96",X"44",X"69",X"9A",X"CD",X"B8",X"43",X"46",X"89",X"9B",X"DE",X"B7",X"32",
		X"35",X"89",X"99",X"AD",X"FF",X"DB",X"97",X"67",X"87",X"53",X"33",X"33",X"46",X"50",X"00",X"6D",
		X"FC",X"7F",X"FF",X"F5",X"00",X"28",X"C9",X"9F",X"FF",X"71",X"01",X"AC",X"38",X"FF",X"F0",X"00",
		X"AE",X"75",X"FF",X"E0",X"00",X"7D",X"76",X"FF",X"F2",X"00",X"7F",X"D6",X"FF",X"F4",X"00",X"6C",
		X"99",X"FF",X"71",X"00",X"99",X"5E",X"FF",X"20",X"08",X"C5",X"8F",X"F8",X"00",X"4D",X"86",X"FF",
		X"90",X"00",X"C7",X"6F",X"FC",X"00",X"0C",X"87",X"FF",X"60",X"05",X"C5",X"BF",X"F0",X"00",X"B9",
		X"6F",X"FD",X"00",X"4F",X"78",X"FF",X"10",X"0C",X"9A",X"FF",X"40",X"09",X"B9",X"FF",X"B0",X"07",
		X"C8",X"DF",X"F0",X"04",X"E9",X"EF",X"F0",X"03",X"E6",X"FF",X"F0",X"08",X"F5",X"FF",X"F0",X"0D",
		X"E5",X"FF",X"F0",X"0F",X"95",X"FF",X"50",X"0F",X"30",X"FF",X"00",X"4F",X"03",X"FF",X"00",X"FF",
		X"0D",X"FF",X"00",X"F6",X"0F",X"FF",X"04",X"F0",X"0F",X"FC",X"0F",X"F0",X"4F",X"FD",X"0D",X"81",
		X"FF",X"FC",X"04",X"90",X"FF",X"EC",X"00",X"E0",X"CF",X"F4",X"00",X"20",X"FF",X"F3",X"00",X"02",
		X"EF",X"F5",X"09",X"05",X"FF",X"F6",X"0C",X"00",X"FF",X"F6",X"0C",X"09",X"9F",X"FB",X"0C",X"00",
		X"9F",X"F6",X"0F",X"0F",X"1F",X"F8",X"0A",X"0F",X"0F",X"F7",X"36",X"0F",X"0F",X"F7",X"81",X"0F",
		X"0F",X"F4",X"40",X"0F",X"0F",X"F7",X"90",X"0F",X"0F",X"EF",X"10",X"0F",X"0F",X"FF",X"00",X"0F",
		X"0F",X"FF",X"0F",X"0F",X"0F",X"FF",X"00",X"0F",X"0F",X"FF",X"0F",X"0F",X"0F",X"FF",X"0B",X"0F",
		X"0F",X"FF",X"00",X"0F",X"0F",X"F7",X"0F",X"0F",X"0F",X"F0",X"A0",X"07",X"7F",X"F0",X"F0",X"50",
		X"F8",X"F0",X"F0",X"81",X"FF",X"F0",X"F0",X"F0",X"FE",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"F0",
		X"FD",X"F0",X"F0",X"F0",X"FF",X"F0",X"81",X"C1",X"FF",X"FC",X"00",X"0F",X"FF",X"F9",X"00",X"0F",
		X"FF",X"3F",X"03",X"0F",X"FF",X"E4",X"00",X"0F",X"9F",X"6D",X"06",X"0D",X"FF",X"F0",X"50",X"4D",
		X"DF",X"07",X"0F",X"0A",X"5F",X"F0",X"F0",X"F0",X"FF",X"F0",X"F0",X"0E",X"0F",X"FF",X"00",X"00",
		X"FF",X"F0",X"F0",X"B0",X"8F",X"FD",X"B0",X"00",X"FF",X"FF",X"F0",X"B0",X"FF",X"FF",X"F0",X"71",
		X"FF",X"F0",X"F0",X"B0",X"FF",X"FF",X"00",X"01",X"F1",X"F5",X"F0",X"F0",X"9E",X"1F",X"F9",X"0F",
		X"0F",X"FF",X"30",X"B0",X"FF",X"AF",X"9F",X"01",X"0F",X"F0",X"F0",X"F0",X"FD",X"F0",X"F0",X"F9",
		X"0F",X"F0",X"F0",X"F0",X"FF",X"FF",X"08",X"0F",X"FF",X"0F",X"00",X"F0",X"FF",X"EF",X"0F",X"0D",
		X"FB",X"F0",X"F0",X"FF",X"F4",X"F0",X"00",X"FF",X"F8",X"0B",X"0F",X"CF",X"06",X"F0",X"FE",X"9F",
		X"F2",X"0F",X"0F",X"F0",X"F0",X"CF",X"DF",X"0F",X"0B",X"F4",X"8F",X"FE",X"0F",X"0F",X"F0",X"20",
		X"0F",X"3F",X"00",X"F0",X"3E",X"FF",X"0F",X"00",X"F0",X"0F",X"0B",X"9F",X"F0",X"08",X"0F",X"0F",
		X"FF",X"30",X"F0",X"FF",X"00",X"60",X"FF",X"0A",X"FC",X"0F",X"0F",X"FF",X"0F",X"5F",X"50",X"FF",
		X"00",X"F0",X"F7",X"0F",X"6F",X"40",X"FF",X"0A",X"F0",X"F0",X"0F",X"0F",X"F0",X"FF",X"0F",X"30",
		X"F0",X"0F",X"04",X"F0",X"8F",X"0F",X"F0",X"F7",X"0F",X"B0",X"F0",X"0F",X"00",X"F2",X"0F",X"05",
		X"F0",X"0F",X"00",X"F0",X"0F",X"00",X"FF",X"0F",X"F0",X"FF",X"0D",X"F0",X"3F",X"0F",X"F0",X"FF",
		X"81",X"FF",X"03",X"F0",X"0F",X"F0",X"FF",X"0F",X"F0",X"0F",X"E0",X"0F",X"00",X"F7",X"05",X"F3",
		X"0F",X"F0",X"FF",X"00",X"FF",X"00",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"FF",X"09",X"F8",
		X"0F",X"F7",X"0D",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"F0",X"0F",X"C0",X"0F",X"D0",X"FF",X"81",
		X"7F",X"E0",X"0F",X"B0",X"5F",X"90",X"FF",X"00",X"DF",X"00",X"FF",X"F0",X"FF",X"00",X"FF",X"00",
		X"FF",X"24",X"FB",X"04",X"FE",X"30",X"CF",X"06",X"F8",X"05",X"FF",X"91",X"FF",X"0F",X"F0",X"0F",
		X"F0",X"FF",X"F9",X"0F",X"E0",X"FF",X"00",X"FF",X"90",X"FF",X"00",X"F6",X"0F",X"F0",X"0F",X"D0",
		X"FF",X"00",X"F0",X"0F",X"F0",X"0F",X"0F",X"F0",X"0F",X"B0",X"FF",X"1F",X"00",X"F1",X"0F",X"F5",
		X"F0",X"0F",X"40",X"FF",X"FF",X"09",X"F0",X"65",X"00",X"00",X"00",X"CD",X"0F",X"FB",X"FF",X"0F",
		X"00",X"A3",X"90",X"03",X"50",X"00",X"CF",X"C0",X"0E",X"EB",X"00",X"FF",X"8F",X"FF",X"3C",X"FF",
		X"00",X"FF",X"00",X"FC",X"0F",X"F0",X"0F",X"CC",X"FD",X"08",X"E9",X"FB",X"02",X"C6",X"00",X"99",
		X"17",X"F4",X"01",X"D1",X"7E",X"EF",X"F0",X"7B",X"26",X"E9",X"FB",X"36",X"73",X"87",X"59",X"A5",
		X"89",X"CC",X"47",X"DA",X"9C",X"98",X"96",X"69",X"86",X"89",X"97",X"89",X"98",X"AB",X"AA",X"79",
		X"87",X"98",X"78",X"A9",X"99",X"89",X"88",X"99",X"98",X"68",X"87",X"79",X"88",X"88",X"70",X"70",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70",
		X"88",X"89",X"89",X"99",X"87",X"67",X"89",X"AA",X"98",X"76",X"67",X"9A",X"98",X"76",X"78",X"AB",
		X"97",X"67",X"AB",X"97",X"79",X"BA",X"64",X"8B",X"86",X"7B",X"A3",X"5C",X"B5",X"4D",X"93",X"8F",
		X"66",X"E8",X"1A",X"81",X"7B",X"3C",X"F6",X"DF",X"6B",X"E2",X"77",X"06",X"50",X"98",X"7F",X"8C",
		X"F6",X"E9",X"0C",X"03",X"90",X"BA",X"9F",X"7D",X"F3",X"E4",X"59",X"08",X"35",X"F6",X"DF",X"4F",
		X"46",X"81",X"B0",X"9C",X"5F",X"5F",X"A9",X"91",X"B0",X"B1",X"BA",X"9D",X"7E",X"3C",X"09",X"0C",
		X"3F",X"6F",X"5E",X"1B",X"0B",X"3E",X"6D",X"7A",X"64",X"91",X"B5",X"F5",X"F3",X"B2",X"65",X"5C",
		X"7F",X"5E",X"27",X"56",X"B7",X"F4",X"E4",X"85",X"3C",X"4F",X"5E",X"59",X"74",X"93",X"E6",X"E8",
		X"99",X"1A",X"2D",X"6C",X"B7",X"A1",X"94",X"9B",X"7E",X"5A",X"83",X"94",X"CB",X"9D",X"48",X"62",
		X"C8",X"BE",X"48",X"53",X"C6",X"9D",X"48",X"82",X"A5",X"7F",X"79",X"B1",X"4B",X"6B",X"E5",X"6B",
		X"44",X"E9",X"6C",X"A3",X"6B",X"79",X"C8",X"26",X"B8",X"9D",X"93",X"6B",X"75",X"DC",X"44",X"9A",
		X"4C",X"E7",X"47",X"A8",X"7C",X"94",X"59",X"C7",X"8B",X"94",X"4A",X"D9",X"79",X"77",X"8A",X"BA",
		X"64",X"4C",X"F5",X"37",X"B7",X"99",X"89",X"57",X"A7",X"98",X"6B",X"A6",X"47",X"B3",X"EF",X"82",
		X"B6",X"78",X"99",X"89",X"88",X"87",X"88",X"78",X"78",X"88",X"88",X"98",X"88",X"88",X"88",X"89",
		X"87",X"78",X"98",X"87",X"88",X"97",X"78",X"89",X"98",X"89",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"98",X"89",X"88",X"88",X"88",X"88",
		X"88",X"98",X"98",X"88",X"98",X"88",X"88",X"88",X"98",X"79",X"88",X"78",X"88",X"88",X"88",X"70",
		X"88",X"88",X"98",X"89",X"88",X"88",X"88",X"88",X"79",X"88",X"98",X"89",X"78",X"88",X"78",X"78",
		X"88",X"88",X"89",X"88",X"88",X"87",X"88",X"89",X"89",X"98",X"98",X"89",X"78",X"78",X"87",X"98",
		X"99",X"89",X"88",X"87",X"87",X"98",X"99",X"8A",X"78",X"87",X"87",X"97",X"97",X"97",X"97",X"87",
		X"87",X"88",X"89",X"98",X"98",X"97",X"97",X"98",X"98",X"99",X"79",X"79",X"79",X"88",X"97",X"97",
		X"98",X"99",X"89",X"78",X"77",X"97",X"A7",X"98",X"79",X"69",X"88",X"A7",X"97",X"89",X"79",X"79",
		X"97",X"97",X"87",X"89",X"79",X"78",X"87",X"97",X"99",X"88",X"78",X"86",X"98",X"8A",X"78",X"96",
		X"89",X"8A",X"97",X"98",X"7A",X"97",X"A8",X"79",X"77",X"A9",X"89",X"76",X"99",X"89",X"97",X"78",
		X"77",X"99",X"77",X"88",X"78",X"A8",X"77",X"88",X"89",X"97",X"78",X"99",X"89",X"97",X"78",X"A9",
		X"88",X"88",X"78",X"9A",X"77",X"89",X"98",X"78",X"88",X"78",X"99",X"87",X"79",X"A9",X"76",X"88",
		X"99",X"67",X"89",X"89",X"87",X"78",X"99",X"87",X"78",X"99",X"89",X"87",X"99",X"77",X"88",X"70",
		X"88",X"88",X"88",X"88",X"79",X"84",X"99",X"C9",X"59",X"B6",X"5A",X"E8",X"69",X"9C",X"65",X"AB",
		X"93",X"8C",X"75",X"5A",X"B6",X"58",X"BB",X"46",X"CB",X"55",X"9C",X"75",X"5B",X"C6",X"49",X"C9",
		X"48",X"9A",X"75",X"9C",X"95",X"6B",X"C6",X"59",X"BA",X"55",X"9C",X"95",X"7C",X"A6",X"6A",X"B7",
		X"66",X"AC",X"64",X"7C",X"A6",X"59",X"B9",X"55",X"AB",X"74",X"6B",X"C6",X"58",X"CA",X"54",X"9C",
		X"A5",X"59",X"C9",X"55",X"AD",X"95",X"59",X"C9",X"55",X"9C",X"95",X"6A",X"B7",X"57",X"CC",X"74",
		X"7B",X"C7",X"46",X"CC",X"63",X"8D",X"B5",X"37",X"EC",X"43",X"9E",X"B4",X"4A",X"E9",X"34",X"BE",
		X"83",X"4B",X"E7",X"36",X"DD",X"53",X"6E",X"D5",X"28",X"EC",X"43",X"9E",X"A3",X"3A",X"E9",X"34",
		X"AE",X"92",X"5C",X"E7",X"25",X"CD",X"63",X"6C",X"E6",X"36",X"DE",X"62",X"7D",X"D5",X"26",X"DD",
		X"52",X"6D",X"E6",X"25",X"DE",X"72",X"5D",X"E8",X"24",X"BF",X"A2",X"39",X"EB",X"42",X"6D",X"F9",
		X"33",X"8D",X"E6",X"32",X"8E",X"F7",X"22",X"7E",X"F9",X"21",X"7E",X"FB",X"31",X"3B",X"FE",X"62",
		X"26",X"EF",X"C6",X"13",X"7F",X"FB",X"41",X"39",X"FF",X"A4",X"13",X"9F",X"F9",X"52",X"28",X"DF",
		X"D7",X"32",X"4A",X"DF",X"D6",X"32",X"39",X"EE",X"E7",X"31",X"26",X"DF",X"FB",X"63",X"12",X"6D",
		X"FE",X"D6",X"31",X"25",X"AE",X"FE",X"87",X"22",X"26",X"AE",X"EE",X"97",X"33",X"24",X"7B",X"DD",
		X"EB",X"84",X"33",X"35",X"6B",X"DE",X"DB",X"98",X"34",X"23",X"56",X"BB",X"EE",X"EB",X"87",X"34",
		X"32",X"55",X"7C",X"CC",X"ED",X"DB",X"75",X"33",X"33",X"57",X"79",X"DE",X"CD",X"D9",X"99",X"65",
		X"44",X"45",X"66",X"8A",X"BA",X"AB",X"BA",X"89",X"98",X"65",X"66",X"66",X"77",X"88",X"99",X"AA",
		X"99",X"9A",X"98",X"77",X"78",X"77",X"66",X"67",X"89",X"98",X"87",X"89",X"99",X"99",X"99",X"88",
		X"98",X"88",X"87",X"77",X"77",X"77",X"78",X"88",X"88",X"88",X"89",X"89",X"89",X"89",X"89",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"78",X"88",X"88",X"88",X"88",X"88",X"98",X"98",X"88",
		X"98",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"98",X"88",X"77",X"88",X"88",X"87",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"70",
		X"86",X"66",X"78",X"99",X"98",X"77",X"89",X"BB",X"B9",X"75",X"55",X"68",X"99",X"97",X"76",X"8A",
		X"BC",X"B9",X"65",X"44",X"68",X"AA",X"98",X"66",X"79",X"BC",X"CB",X"95",X"33",X"47",X"9A",X"B9",
		X"76",X"68",X"AC",X"DD",X"B7",X"43",X"34",X"69",X"AA",X"96",X"56",X"9C",X"DD",X"C9",X"64",X"23",
		X"57",X"9A",X"A8",X"66",X"8A",X"CC",X"CB",X"97",X"33",X"35",X"79",X"AA",X"97",X"89",X"AB",X"9A",
		X"98",X"65",X"45",X"67",X"89",X"98",X"98",X"99",X"99",X"99",X"88",X"77",X"77",X"78",X"89",X"99",
		X"99",X"89",X"98",X"88",X"77",X"77",X"77",X"88",X"99",X"99",X"88",X"89",X"98",X"88",X"77",X"67",
		X"88",X"89",X"99",X"98",X"88",X"87",X"88",X"88",X"77",X"77",X"88",X"88",X"89",X"88",X"98",X"88",
		X"88",X"88",X"78",X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"88",X"88",X"88",X"88",X"89",X"88",
		X"87",X"78",X"88",X"88",X"98",X"78",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"89",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"78",X"88",X"88",X"88",X"89",X"87",
		X"88",X"88",X"78",X"89",X"98",X"98",X"89",X"88",X"99",X"88",X"88",X"79",X"97",X"97",X"77",X"64",
		X"35",X"9C",X"FC",X"40",X"05",X"64",X"AF",X"FF",X"60",X"0A",X"E7",X"0A",X"FF",X"81",X"08",X"F9",
		X"01",X"FF",X"F0",X"08",X"FE",X"00",X"FF",X"F0",X"0B",X"FC",X"00",X"FF",X"F0",X"06",X"FC",X"00",
		X"FF",X"F0",X"01",X"FF",X"00",X"FF",X"F0",X"08",X"FF",X"00",X"FF",X"F0",X"0D",X"FC",X"00",X"FF",
		X"F0",X"0D",X"F0",X"02",X"FF",X"50",X"0F",X"F0",X"09",X"FF",X"B0",X"9F",X"B0",X"0F",X"FF",X"00",
		X"FF",X"00",X"7F",X"F3",X"03",X"FB",X"00",X"FF",X"F0",X"0F",X"F0",X"0A",X"FF",X"60",X"CF",X"30",
		X"4F",X"FF",X"00",X"FC",X"00",X"FF",X"F0",X"0F",X"F0",X"0C",X"FF",X"71",X"FF",X"00",X"9F",X"F6",
		X"0E",X"F0",X"07",X"FF",X"60",X"EF",X"00",X"8F",X"F8",X"0F",X"F0",X"09",X"FF",X"E0",X"FF",X"00",
		X"AF",X"F0",X"0F",X"F0",X"09",X"FF",X"00",X"FC",X"01",X"FF",X"A0",X"8F",X"00",X"CF",X"FB",X"0F",
		X"F0",X"0A",X"FF",X"00",X"F9",X"0B",X"AF",X"90",X"0F",X"00",X"F7",X"FF",X"0F",X"F0",X"1D",X"3F",
		X"F0",X"FF",X"02",X"B3",X"FF",X"0F",X"F0",X"5E",X"0F",X"F0",X"FF",X"01",X"F0",X"FF",X"00",X"F1",
		X"0F",X"71",X"FF",X"0F",X"F0",X"4F",X"00",X"F7",X"0F",X"F0",X"CF",X"00",X"FF",X"0E",X"F0",X"6F",
		X"25",X"F9",X"CE",X"7E",X"B3",X"6D",X"55",X"97",X"9B",X"85",X"5A",X"68",X"B7",X"7A",X"86",X"98",
		X"4A",X"C2",X"5D",X"85",X"BB",X"68",X"96",X"99",X"68",X"86",X"9B",X"77",X"97",X"79",X"78",X"A9",
		X"78",X"98",X"78",X"98",X"98",X"79",X"87",X"89",X"87",X"88",X"88",X"88",X"99",X"88",X"89",X"88",
		X"88",X"89",X"89",X"88",X"89",X"88",X"88",X"78",X"98",X"89",X"88",X"88",X"79",X"89",X"98",X"78",
		X"87",X"89",X"88",X"98",X"89",X"87",X"89",X"88",X"89",X"88",X"88",X"99",X"78",X"98",X"78",X"89",
		X"88",X"89",X"77",X"89",X"97",X"89",X"97",X"78",X"98",X"78",X"98",X"88",X"89",X"87",X"99",X"88",
		X"88",X"88",X"88",X"98",X"88",X"88",X"98",X"88",X"87",X"88",X"89",X"88",X"88",X"88",X"70",X"70",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70",
		X"88",X"89",X"88",X"88",X"88",X"88",X"89",X"A8",X"54",X"8C",X"EC",X"63",X"36",X"9B",X"CC",X"B9",
		X"53",X"37",X"CE",X"C7",X"44",X"8B",X"CA",X"75",X"48",X"CB",X"53",X"2B",X"EF",X"E8",X"31",X"12",
		X"8E",X"FF",X"C4",X"00",X"7D",X"FF",X"63",X"35",X"78",X"AE",X"EE",X"93",X"10",X"5C",X"EE",X"C7",
		X"43",X"33",X"8E",X"FF",X"E6",X"10",X"06",X"CF",X"FD",X"63",X"22",X"5C",X"FF",X"F8",X"40",X"06",
		X"CF",X"FB",X"62",X"23",X"7C",X"FF",X"D6",X"20",X"29",X"DF",X"E9",X"43",X"34",X"9D",X"FE",X"B4",
		X"11",X"4A",X"CE",X"C7",X"33",X"49",X"CD",X"D9",X"43",X"36",X"BD",X"DB",X"64",X"35",X"AC",X"DB",
		X"74",X"46",X"9B",X"B9",X"76",X"67",X"9A",X"AA",X"86",X"66",X"8A",X"BA",X"86",X"57",X"9B",X"B9",
		X"76",X"67",X"89",X"BA",X"97",X"55",X"79",X"BB",X"96",X"67",X"89",X"99",X"99",X"87",X"77",X"89",
		X"99",X"77",X"78",X"88",X"89",X"99",X"97",X"76",X"79",X"9A",X"98",X"77",X"77",X"89",X"99",X"98",
		X"77",X"78",X"99",X"99",X"87",X"77",X"89",X"A9",X"97",X"77",X"89",X"99",X"98",X"77",X"78",X"99",
		X"98",X"77",X"78",X"89",X"88",X"88",X"88",X"88",X"99",X"87",X"77",X"89",X"99",X"98",X"77",X"78",
		X"99",X"99",X"87",X"77",X"89",X"99",X"87",X"78",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"77",
		X"88",X"88",X"88",X"88",X"87",X"88",X"99",X"87",X"77",X"88",X"99",X"88",X"88",X"87",X"88",X"99",
		X"88",X"88",X"98",X"88",X"88",X"98",X"87",X"88",X"99",X"88",X"78",X"88",X"88",X"88",X"88",X"78",
		X"99",X"98",X"87",X"88",X"89",X"88",X"88",X"88",X"99",X"88",X"88",X"88",X"99",X"98",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"87",X"88",X"99",X"88",X"88",X"88",X"99",X"98",X"87",X"70",
		X"88",X"98",X"88",X"98",X"88",X"97",X"96",X"C2",X"C7",X"89",X"98",X"78",X"88",X"88",X"78",X"88",
		X"88",X"89",X"79",X"D5",X"5C",X"87",X"5A",X"96",X"86",X"EC",X"65",X"B6",X"79",X"89",X"6D",X"A5",
		X"A1",X"5D",X"3C",X"7D",X"76",X"7C",X"0C",X"5C",X"2C",X"8B",X"94",X"A5",X"67",X"F8",X"89",X"08",
		X"F3",X"8A",X"A3",X"6E",X"89",X"93",X"A8",X"5B",X"D3",X"B8",X"46",X"8B",X"D2",X"B4",X"98",X"D7",
		X"96",X"74",X"F4",X"5C",X"A4",X"7B",X"C9",X"71",X"4D",X"D3",X"C8",X"37",X"A5",X"7F",X"96",X"81",
		X"9F",X"5B",X"36",X"9D",X"3A",X"B5",X"2F",X"A2",X"FA",X"37",X"A4",X"E5",X"7C",X"76",X"3D",X"8A",
		X"B6",X"46",X"DA",X"58",X"79",X"96",X"9B",X"28",X"E4",X"C9",X"66",X"B0",X"B8",X"C6",X"58",X"97",
		X"B7",X"7D",X"56",X"C6",X"8C",X"73",X"6D",X"E4",X"86",X"92",X"F6",X"BA",X"54",X"B7",X"89",X"A7",
		X"A6",X"92",X"D7",X"D5",X"63",X"F9",X"93",X"68",X"AC",X"C6",X"16",X"AC",X"6C",X"C4",X"39",X"6F",
		X"69",X"1F",X"5B",X"3C",X"87",X"C5",X"3D",X"5D",X"95",X"1F",X"2C",X"8B",X"55",X"6E",X"78",X"97",
		X"77",X"9B",X"84",X"99",X"7A",X"66",X"97",X"A7",X"95",X"D6",X"B5",X"98",X"79",X"9A",X"28",X"6E",
		X"C3",X"67",X"E7",X"89",X"84",X"A9",X"A7",X"96",X"84",X"AB",X"B4",X"8A",X"76",X"99",X"AC",X"66",
		X"66",X"B9",X"96",X"87",X"AA",X"83",X"98",X"9A",X"C6",X"39",X"87",X"BD",X"58",X"59",X"C2",X"B8",
		X"D3",X"A6",X"A6",X"8B",X"85",X"88",X"A9",X"58",X"86",X"9C",X"89",X"35",X"C8",X"79",X"B8",X"65",
		X"BC",X"38",X"BC",X"65",X"7C",X"49",X"9A",X"69",X"79",X"93",X"B7",X"B8",X"9A",X"75",X"8C",X"87",
		X"96",X"89",X"89",X"77",X"5E",X"B6",X"2A",X"A6",X"99",X"87",X"97",X"87",X"8C",X"77",X"6A",X"68",
		X"7B",X"87",X"6A",X"89",X"A5",X"6D",X"94",X"8C",X"B6",X"66",X"7C",X"AB",X"3B",X"49",X"98",X"B9",
		X"75",X"87",X"DA",X"85",X"6A",X"B4",X"8B",X"48",X"B6",X"96",X"C8",X"57",X"B8",X"98",X"7B",X"65",
		X"9B",X"9B",X"47",X"99",X"7A",X"88",X"69",X"97",X"87",X"89",X"88",X"97",X"6B",X"78",X"7B",X"87",
		X"6B",X"67",X"9A",X"97",X"67",X"99",X"95",X"A8",X"89",X"87",X"88",X"7B",X"79",X"68",X"77",X"A7",
		X"79",X"A7",X"86",X"6A",X"A9",X"95",X"79",X"89",X"98",X"6A",X"79",X"78",X"99",X"78",X"9A",X"57",
		X"B8",X"6B",X"77",X"C7",X"66",X"A7",X"A9",X"95",X"7A",X"6A",X"88",X"98",X"6A",X"96",X"8B",X"97",
		X"88",X"88",X"99",X"88",X"97",X"97",X"86",X"7A",X"C7",X"79",X"59",X"A8",X"8A",X"58",X"A8",X"A7",
		X"75",X"CB",X"57",X"8A",X"69",X"88",X"8A",X"78",X"77",X"A9",X"78",X"68",X"99",X"68",X"A8",X"68",
		X"B8",X"57",X"99",X"A8",X"76",X"89",X"C6",X"5B",X"88",X"6A",X"79",X"79",X"7A",X"94",X"A8",X"97",
		X"B4",X"98",X"98",X"96",X"9A",X"77",X"89",X"78",X"89",X"6A",X"99",X"76",X"89",X"89",X"A6",X"97",
		X"89",X"A6",X"89",X"8A",X"69",X"69",X"99",X"79",X"68",X"A7",X"79",X"96",X"A9",X"86",X"79",X"99",
		X"97",X"78",X"99",X"79",X"88",X"98",X"88",X"78",X"B8",X"87",X"97",X"98",X"97",X"99",X"79",X"96",
		X"79",X"B9",X"77",X"96",X"8A",X"87",X"89",X"97",X"78",X"97",X"A8",X"96",X"6A",X"87",X"99",X"79",
		X"97",X"88",X"88",X"8B",X"76",X"8A",X"79",X"88",X"87",X"99",X"77",X"99",X"88",X"88",X"69",X"70",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",
		X"88",X"99",X"89",X"88",X"78",X"88",X"89",X"A9",X"B7",X"5A",X"57",X"86",X"98",X"9B",X"BA",X"3C",
		X"48",X"85",X"87",X"AB",X"CC",X"0F",X"27",X"93",X"A6",X"9A",X"CD",X"64",X"95",X"96",X"67",X"8A",
		X"BE",X"C0",X"F1",X"7A",X"29",X"6B",X"AE",X"E0",X"F0",X"6B",X"1C",X"4A",X"BE",X"F0",X"F0",X"6B",
		X"0B",X"58",X"BD",X"F0",X"F3",X"6B",X"1B",X"59",X"CD",X"F0",X"A6",X"5B",X"27",X"69",X"DB",X"F0",
		X"B6",X"3C",X"07",X"79",X"EC",X"F0",X"F3",X"3E",X"09",X"69",X"EE",X"F0",X"F1",X"1E",X"09",X"5B",
		X"DF",X"F0",X"F1",X"2C",X"19",X"4F",X"DF",X"0F",X"50",X"F0",X"87",X"9F",X"FF",X"0F",X"24",X"93",
		X"B3",X"FE",X"F0",X"F6",X"0E",X"28",X"6B",X"FF",X"0F",X"71",X"D1",X"66",X"CF",X"F3",X"B9",X"0D",
		X"07",X"88",X"FF",X"59",X"81",X"B4",X"4A",X"9F",X"F3",X"AA",X"0B",X"53",X"8B",X"FF",X"0B",X"D0",
		X"97",X"39",X"CF",X"F0",X"9F",X"06",X"A4",X"7E",X"FE",X"07",X"E0",X"2A",X"77",X"FF",X"92",X"6A",
		X"64",X"67",X"8A",X"ED",X"73",X"57",X"97",X"79",X"BE",X"C7",X"43",X"78",X"77",X"9A",X"DC",X"63",
		X"37",X"97",X"89",X"BD",X"B6",X"34",X"69",X"88",X"9C",X"DA",X"44",X"56",X"98",X"AC",X"F9",X"23",
		X"88",X"46",X"9E",X"FF",X"10",X"C6",X"09",X"97",X"FF",X"00",X"F6",X"09",X"A5",X"FF",X"71",X"C8",
		X"08",X"B4",X"DF",X"F0",X"4D",X"13",X"94",X"9F",X"F7",X"0E",X"60",X"88",X"6D",X"FF",X"05",X"D0",
		X"59",X"39",X"FF",X"60",X"E5",X"08",X"65",X"FF",X"F0",X"7C",X"06",X"A4",X"8F",X"F6",X"0E",X"60",
		X"77",X"6E",X"FF",X"06",X"C0",X"3A",X"68",X"FF",X"81",X"D8",X"05",X"85",X"BF",X"F0",X"2D",X"21",
		X"97",X"7F",X"FB",X"0C",X"B0",X"3A",X"59",X"FF",X"00",X"E3",X"09",X"96",X"FF",X"B0",X"CD",X"02",
		X"C6",X"9F",X"F0",X"2E",X"30",X"89",X"5F",X"F7",X"0B",X"D0",X"3D",X"6A",X"FF",X"02",X"E5",X"07",
		X"A4",X"EF",X"71",X"AE",X"03",X"D7",X"BF",X"F0",X"3F",X"40",X"AA",X"5F",X"F3",X"0B",X"B0",X"2C",
		X"7B",X"FF",X"04",X"F4",X"0B",X"B7",X"FF",X"20",X"DA",X"02",X"C6",X"CF",X"D0",X"5F",X"30",X"BA",
		X"9F",X"F2",X"0E",X"81",X"5B",X"6D",X"F7",X"07",X"D0",X"0C",X"9B",X"FF",X"01",X"F8",X"07",X"B7",
		X"EF",X"50",X"8C",X"01",X"B9",X"BF",X"F0",X"3F",X"71",X"9B",X"8F",X"F3",X"0B",X"B0",X"2C",X"7B",
		X"FC",X"04",X"F4",X"0A",X"A9",X"FF",X"40",X"CA",X"03",X"B7",X"CF",X"90",X"6F",X"20",X"BA",X"BF",
		X"F2",X"1F",X"81",X"6C",X"6E",X"F6",X"07",X"E0",X"0C",X"9B",X"FF",X"02",X"F7",X"07",X"B7",X"FF",
		X"40",X"9C",X"01",X"C8",X"CF",X"F0",X"4F",X"50",X"9A",X"8F",X"F3",X"0B",X"B0",X"2B",X"7C",X"FC",
		X"04",X"F3",X"0A",X"AA",X"FF",X"20",X"D9",X"05",X"B7",X"DF",X"A0",X"4F",X"20",X"AA",X"BF",X"F1",
		X"0D",X"90",X"5B",X"8E",X"F6",X"06",X"E1",X"0B",X"9B",X"FF",X"20",X"D8",X"05",X"A8",X"EF",X"60",
		X"7D",X"00",X"B9",X"CF",X"F0",X"1D",X"90",X"6B",X"8F",X"F6",X"07",X"C0",X"0B",X"9C",X"FF",X"01",
		X"E7",X"07",X"B9",X"FF",X"40",X"9D",X"00",X"B9",X"CF",X"F0",X"2F",X"71",X"7B",X"9F",X"F6",X"08",
		X"C0",X"0B",X"9C",X"FF",X"02",X"F7",X"07",X"B9",X"FF",X"50",X"9C",X"00",X"B9",X"AF",X"F0",X"1F",
		X"90",X"6B",X"8F",X"F5",X"06",X"E0",X"0B",X"9C",X"FF",X"12",X"F9",X"06",X"B8",X"EF",X"40",X"7E",
		X"00",X"B9",X"BF",X"D0",X"3F",X"40",X"8A",X"BF",X"F4",X"0C",X"B0",X"5B",X"8D",X"F7",X"04",X"E1",
		X"09",X"BC",X"FF",X"20",X"DA",X"04",X"C8",X"EF",X"60",X"6E",X"00",X"AA",X"CF",X"F0",X"1F",X"81",
		X"6C",X"BF",X"F4",X"0B",X"C0",X"0B",X"9D",X"F7",X"05",X"E1",X"09",X"BC",X"FF",X"01",X"E8",X"06",
		X"BB",X"FF",X"50",X"BB",X"01",X"BA",X"EF",X"71",X"6D",X"10",X"8A",X"CF",X"C0",X"2E",X"60",X"7B",
		X"CF",X"F3",X"0C",X"B0",X"3B",X"9F",X"F6",X"09",X"C0",X"2B",X"9D",X"F7",X"07",X"C0",X"09",X"AD",
		X"F9",X"03",X"D3",X"08",X"BD",X"FC",X"03",X"E5",X"08",X"BC",X"FF",X"01",X"EA",X"06",X"DB",X"FF",
		X"40",X"DB",X"03",X"BA",X"FF",X"50",X"9C",X"00",X"99",X"DF",X"71",X"4F",X"30",X"9B",X"DF",X"D0",
		X"1F",X"81",X"7C",X"CF",X"F2",X"0D",X"A0",X"5B",X"CF",X"F4",X"0D",X"B0",X"6C",X"BF",X"F4",X"0C",
		X"C0",X"4B",X"9F",X"F6",X"09",X"C0",X"0A",X"AC",X"F6",X"06",X"D1",X"09",X"BD",X"F9",X"03",X"F4",
		X"09",X"CD",X"FC",X"00",X"E8",X"07",X"CC",X"FF",X"30",X"CC",X"03",X"BB",X"FF",X"60",X"AC",X"01",
		X"B9",X"DF",X"60",X"6D",X"00",X"9B",X"DF",X"90",X"2E",X"50",X"7C",X"DF",X"F2",X"1C",X"B0",X"5B",
		X"BF",X"F6",X"0B",X"C0",X"2B",X"AD",X"F6",X"07",X"C0",X"09",X"9C",X"F8",X"03",X"D4",X"08",X"BC",
		X"FF",X"01",X"D8",X"07",X"BB",X"FF",X"50",X"AA",X"03",X"BA",X"EF",X"71",X"9C",X"00",X"99",X"CF",
		X"90",X"4C",X"30",X"9B",X"DF",X"D0",X"1E",X"60",X"7C",X"DF",X"F4",X"1D",X"B0",X"5C",X"AF",X"F6",
		X"09",X"C0",X"1A",X"9C",X"F8",X"03",X"D3",X"08",X"BD",X"FF",X"01",X"D7",X"06",X"BB",X"FF",X"60",
		X"CB",X"04",X"BA",X"EF",X"60",X"8C",X"00",X"A9",X"CF",X"B0",X"1D",X"50",X"7B",X"DF",X"F3",X"0C",
		X"B0",X"5B",X"AF",X"F7",X"08",X"C0",X"09",X"9C",X"F9",X"01",X"D5",X"07",X"BD",X"FF",X"20",X"CA",
		X"06",X"BA",X"FF",X"71",X"9C",X"00",X"99",X"DF",X"81",X"2C",X"30",X"7A",X"CF",X"F1",X"0C",X"A0",
		X"6B",X"BF",X"F7",X"08",X"B1",X"29",X"9C",X"F8",X"03",X"B4",X"17",X"AC",X"FE",X"01",X"B8",X"06",
		X"AB",X"FF",X"71",X"9B",X"03",X"99",X"DF",X"81",X"4B",X"31",X"79",X"CF",X"F1",X"1B",X"81",X"6A",
		X"BF",X"F7",X"09",X"B1",X"29",X"AD",X"F8",X"03",X"C4",X"08",X"AD",X"FF",X"21",X"BA",X"16",X"AA",
		X"EF",X"71",X"7B",X"22",X"99",X"CF",X"90",X"3B",X"51",X"7A",X"CF",X"F3",X"1B",X"91",X"6B",X"BF",
		X"F7",X"09",X"B1",X"39",X"9B",X"F9",X"03",X"B5",X"17",X"AC",X"FE",X"12",X"B8",X"17",X"BC",X"FF",
		X"50",X"9A",X"14",X"AA",X"EF",X"60",X"5B",X"10",X"9A",X"DF",X"C0",X"1D",X"71",X"7B",X"DF",X"F4",
		X"0B",X"A0",X"4B",X"AE",X"F7",X"06",X"B2",X"19",X"AD",X"FB",X"02",X"C6",X"07",X"AC",X"FF",X"41",
		X"AA",X"14",X"AA",X"EF",X"71",X"5B",X"21",X"9A",X"DF",X"D0",X"2C",X"71",X"7B",X"CF",X"F4",X"0A",
		X"A0",X"4A",X"9D",X"F8",X"03",X"B4",X"08",X"AC",X"FF",X"31",X"B9",X"16",X"BB",X"FF",X"60",X"8A",
		X"23",X"99",X"CF",X"90",X"4B",X"41",X"8A",X"CF",X"F2",X"2C",X"90",X"6B",X"BF",X"F6",X"08",X"B0",
		X"2A",X"9C",X"F9",X"02",X"C5",X"18",X"AC",X"FF",X"52",X"A9",X"15",X"AA",X"EF",X"60",X"6B",X"12",
		X"A9",X"DF",X"C0",X"2C",X"60",X"7B",X"BF",X"F6",X"1A",X"A1",X"3A",X"9C",X"F8",X"04",X"B3",X"19",
		X"AC",X"FF",X"22",X"B8",X"06",X"AB",X"FF",X"60",X"7B",X"11",X"99",X"CF",X"C0",X"1C",X"61",X"7A",
		X"BF",X"F5",X"19",X"A1",X"39",X"9C",X"F9",X"03",X"B4",X"18",X"AB",X"FF",X"52",X"A9",X"15",X"AA",
		X"EF",X"60",X"6B",X"31",X"89",X"CF",X"F2",X"2B",X"81",X"6A",X"AE",X"F6",X"06",X"A2",X"18",X"9C",
		X"FE",X"33",X"A7",X"26",X"AB",X"EF",X"60",X"7B",X"21",X"89",X"CF",X"D0",X"2B",X"72",X"6A",X"BF",
		X"F6",X"07",X"A2",X"39",X"9C",X"FA",X"03",X"A6",X"27",X"9B",X"FF",X"62",X"99",X"25",X"9A",X"CF",
		X"92",X"69",X"64",X"89",X"BE",X"C4",X"49",X"84",X"79",X"AD",X"F7",X"27",X"94",X"49",X"9C",X"FA",
		X"14",X"A6",X"38",X"9B",X"EE",X"63",X"99",X"35",X"9A",X"DF",X"71",X"5A",X"33",X"89",X"CF",X"C0",
		X"3B",X"82",X"7B",X"BF",X"F6",X"18",X"93",X"49",X"9C",X"FA",X"03",X"B6",X"38",X"AC",X"FF",X"42",
		X"99",X"35",X"9A",X"DF",X"71",X"6A",X"43",X"99",X"CF",X"C1",X"3B",X"72",X"7A",X"BF",X"F6",X"28",
		X"93",X"69",X"9C",X"F8",X"16",X"A5",X"39",X"AC",X"FC",X"23",X"B7",X"27",X"AB",X"EE",X"42",X"99",
		X"36",X"9A",X"CF",X"73",X"79",X"45",X"99",X"BD",X"95",X"69",X"76",X"89",X"99",X"98",X"88",X"87",
		X"89",X"9A",X"B6",X"49",X"94",X"59",X"9B",X"C7",X"67",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"98",X"88",X"88",X"88",X"89",X"98",X"77",X"97",X"68",X"99",X"BB",X"65",X"98",X"57",X"9A",
		X"BC",X"64",X"89",X"46",X"99",X"BE",X"72",X"6A",X"54",X"89",X"BE",X"B3",X"49",X"74",X"79",X"BD",
		X"D4",X"39",X"84",X"69",X"AD",X"E6",X"28",X"A4",X"49",X"9C",X"F9",X"15",X"B6",X"48",X"9B",X"EC",
		X"34",X"98",X"46",X"9A",X"DE",X"53",X"99",X"36",X"99",X"CF",X"71",X"6A",X"54",X"99",X"BF",X"B3",
		X"5A",X"73",X"89",X"BD",X"D5",X"39",X"93",X"69",X"9C",X"F6",X"17",X"A4",X"49",X"9B",X"EB",X"35",
		X"96",X"37",X"9A",X"CD",X"63",X"8A",X"44",X"99",X"BE",X"B4",X"59",X"74",X"79",X"AC",X"E6",X"28",
		X"94",X"59",X"9B",X"EB",X"45",X"A6",X"36",X"99",X"CE",X"73",X"88",X"56",X"99",X"BC",X"95",X"79",
		X"65",X"89",X"AC",X"C6",X"59",X"74",X"89",X"9B",X"D8",X"37",X"96",X"59",X"9A",X"CD",X"64",X"88",
		X"46",X"99",X"BE",X"A3",X"59",X"65",X"89",X"AC",X"D6",X"38",X"84",X"68",X"9B",X"EA",X"46",X"96",
		X"58",X"9A",X"CC",X"75",X"88",X"57",X"99",X"BC",X"95",X"78",X"66",X"89",X"AC",X"B5",X"69",X"75",
		X"79",X"9C",X"C7",X"59",X"85",X"79",X"9B",X"D9",X"47",X"96",X"68",X"9A",X"CC",X"55",X"97",X"57",
		X"99",X"BD",X"83",X"79",X"65",X"99",X"AC",X"C5",X"49",X"84",X"69",X"9B",X"EA",X"46",X"96",X"48",
		X"9A",X"DC",X"54",X"98",X"47",X"99",X"CE",X"93",X"69",X"65",X"99",X"AD",X"C5",X"49",X"74",X"79",
		X"9C",X"E9",X"36",X"95",X"59",X"9B",X"DC",X"44",X"97",X"36",X"99",X"CE",X"83",X"79",X"55",X"99",
		X"BD",X"C4",X"49",X"74",X"79",X"9B",X"E9",X"36",X"96",X"59",X"9B",X"EC",X"44",X"97",X"47",X"99",
		X"DF",X"72",X"79",X"45",X"99",X"BE",X"B4",X"49",X"64",X"79",X"AD",X"E5",X"38",X"84",X"69",X"AC",
		X"F9",X"26",X"94",X"49",X"9B",X"FD",X"43",X"97",X"36",X"9A",X"DF",X"81",X"69",X"55",X"99",X"CF",
		X"C4",X"48",X"74",X"79",X"AD",X"F6",X"07",X"84",X"59",X"9C",X"FB",X"44",X"97",X"47",X"9B",X"DD",
		X"53",X"88",X"46",X"9A",X"CF",X"92",X"69",X"54",X"89",X"BE",X"D3",X"18",X"82",X"59",X"AD",X"F8",
		X"06",X"A4",X"49",X"9C",X"FC",X"24",X"A6",X"37",X"9B",X"FE",X"32",X"97",X"26",X"9A",X"EF",X"81",
		X"6A",X"44",X"99",X"CF",X"D2",X"3A",X"63",X"79",X"AE",X"F5",X"17",X"83",X"69",X"AD",X"F9",X"16",
		X"A4",X"38",X"9C",X"FC",X"34",X"96",X"37",X"9B",X"FF",X"41",X"88",X"36",X"9A",X"DF",X"81",X"69",
		X"45",X"99",X"CF",X"C3",X"49",X"64",X"89",X"BE",X"E4",X"28",X"73",X"69",X"AD",X"F8",X"16",X"94",
		X"59",X"9C",X"FC",X"34",X"95",X"38",X"9B",X"EE",X"42",X"87",X"46",X"9A",X"CE",X"A3",X"69",X"55",
		X"99",X"BE",X"B4",X"49",X"64",X"89",X"BE",X"D4",X"28",X"73",X"69",X"9C",X"F9",X"36",X"95",X"59",
		X"9B",X"EC",X"43",X"87",X"46",X"9A",X"DE",X"83",X"68",X"56",X"99",X"BE",X"B4",X"49",X"74",X"79",
		X"AD",X"E6",X"27",X"84",X"69",X"9B",X"EB",X"44",X"97",X"57",X"9A",X"DD",X"73",X"78",X"56",X"9A",
		X"BE",X"A4",X"69",X"65",X"89",X"AD",X"C5",X"38",X"75",X"79",X"AC",X"D7",X"37",X"85",X"69",X"9B",
		X"D9",X"47",X"96",X"69",X"9B",X"DB",X"45",X"97",X"58",X"9A",X"DB",X"54",X"87",X"58",X"9A",X"CC",
		X"64",X"77",X"57",X"99",X"CC",X"74",X"78",X"57",X"99",X"BC",X"84",X"78",X"67",X"9A",X"BC",X"95",
		X"68",X"66",X"89",X"BC",X"A5",X"58",X"65",X"89",X"AC",X"A6",X"57",X"76",X"89",X"AC",X"B6",X"57",
		X"76",X"79",X"AB",X"B7",X"57",X"76",X"78",X"AB",X"C7",X"57",X"76",X"79",X"AB",X"C8",X"57",X"86",
		X"79",X"AB",X"C8",X"57",X"86",X"79",X"9B",X"C8",X"57",X"86",X"79",X"9B",X"B8",X"57",X"86",X"79",
		X"9B",X"B8",X"57",X"86",X"79",X"9B",X"B8",X"67",X"86",X"79",X"AB",X"B8",X"57",X"87",X"79",X"AB",
		X"B8",X"56",X"77",X"78",X"9B",X"B8",X"66",X"77",X"79",X"9B",X"B8",X"66",X"77",X"79",X"AB",X"B8",
		X"67",X"87",X"89",X"AB",X"B7",X"56",X"77",X"89",X"AB",X"A7",X"56",X"77",X"89",X"AB",X"A7",X"57",
		X"77",X"89",X"AB",X"A7",X"57",X"77",X"89",X"AB",X"A7",X"67",X"77",X"89",X"AB",X"97",X"67",X"77",
		X"89",X"AB",X"97",X"67",X"77",X"89",X"AB",X"97",X"67",X"77",X"89",X"AB",X"96",X"67",X"78",X"99",
		X"AB",X"96",X"67",X"77",X"99",X"AB",X"96",X"67",X"77",X"89",X"AB",X"96",X"67",X"77",X"89",X"AB",
		X"96",X"67",X"77",X"99",X"AB",X"97",X"67",X"77",X"89",X"AB",X"A7",X"67",X"77",X"89",X"AA",X"A7",
		X"67",X"77",X"89",X"9A",X"A8",X"67",X"77",X"89",X"9A",X"A8",X"66",X"77",X"89",X"9A",X"B9",X"66",
		X"77",X"78",X"99",X"A9",X"76",X"77",X"78",X"99",X"A9",X"76",X"78",X"78",X"99",X"AA",X"86",X"78",
		X"78",X"89",X"AA",X"96",X"67",X"77",X"89",X"AA",X"97",X"67",X"77",X"89",X"AA",X"A8",X"67",X"87",
		X"89",X"9A",X"A8",X"67",X"87",X"78",X"9A",X"A9",X"76",X"87",X"78",X"99",X"AA",X"86",X"78",X"78",
		X"89",X"AA",X"86",X"77",X"77",X"89",X"AA",X"86",X"77",X"77",X"89",X"AA",X"97",X"78",X"77",X"89",
		X"AA",X"97",X"76",X"87",X"89",X"AA",X"97",X"67",X"86",X"89",X"9A",X"98",X"67",X"77",X"89",X"9A",
		X"98",X"67",X"87",X"79",X"99",X"99",X"77",X"77",X"78",X"9A",X"A9",X"77",X"78",X"78",X"99",X"A9",
		X"87",X"68",X"78",X"99",X"99",X"87",X"78",X"78",X"89",X"99",X"97",X"77",X"87",X"89",X"99",X"98",
		X"77",X"87",X"89",X"99",X"98",X"77",X"87",X"88",X"99",X"98",X"77",X"77",X"78",X"99",X"98",X"87",
		X"78",X"78",X"89",X"99",X"87",X"78",X"77",X"89",X"99",X"87",X"78",X"77",X"89",X"99",X"98",X"76",
		X"87",X"78",X"99",X"99",X"76",X"87",X"88",X"99",X"99",X"87",X"88",X"78",X"99",X"89",X"88",X"78",
		X"78",X"89",X"89",X"98",X"78",X"78",X"89",X"99",X"88",X"77",X"88",X"88",X"99",X"89",X"87",X"78",
		X"78",X"99",X"99",X"97",X"78",X"78",X"89",X"99",X"88",X"78",X"78",X"88",X"99",X"98",X"77",X"78",
		X"89",X"99",X"98",X"87",X"78",X"88",X"99",X"99",X"88",X"88",X"88",X"99",X"99",X"88",X"70",X"70",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70",
		X"88",X"88",X"87",X"88",X"77",X"78",X"88",X"AF",X"0B",X"0C",X"CF",X"0C",X"FF",X"CF",X"0B",X"C5",
		X"FA",X"90",X"03",X"81",X"71",X"0F",X"08",X"FF",X"93",X"05",X"F6",X"F5",X"AF",X"8E",X"F6",X"FF",
		X"FF",X"AF",X"F6",X"60",X"FF",X"81",X"00",X"9A",X"07",X"01",X"FD",X"A9",X"20",X"00",X"00",X"0F",
		X"0D",X"B2",X"60",X"9F",X"90",X"58",X"F0",X"6F",X"F3",X"07",X"FF",X"9F",X"FF",X"F7",X"FF",X"0F",
		X"FF",X"A0",X"D7",X"F0",X"07",X"A0",X"FB",X"D5",X"07",X"00",X"00",X"04",X"04",X"C0",X"F0",X"FF",
		X"00",X"00",X"B4",X"F9",X"79",X"FF",X"FF",X"FF",X"FF",X"EF",X"2F",X"F7",X"00",X"7F",X"5F",X"FF",
		X"D2",X"04",X"00",X"00",X"D0",X"96",X"00",X"09",X"F6",X"0F",X"F0",X"00",X"60",X"04",X"EF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"EF",X"FF",X"6C",X"B0",X"B9",X"81",X"00",X"00",X"00",
		X"40",X"81",X"00",X"7F",X"D0",X"00",X"40",X"00",X"18",X"FF",X"FE",X"EF",X"FA",X"9F",X"F6",X"5A",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"F1",X"C0",X"00",X"F7",X"20",X"90",X"59",X"30",X"00",X"00",X"00",
		X"00",X"00",X"AF",X"FF",X"E9",X"FA",X"F3",X"9F",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",
		X"00",X"FF",X"19",X"99",X"0A",X"A1",X"30",X"00",X"00",X"00",X"00",X"F0",X"CD",X"53",X"0F",X"A3",
		X"53",X"DA",X"FF",X"FF",X"FF",X"F2",X"FB",X"FF",X"04",X"0F",X"FF",X"0F",X"FF",X"FD",X"90",X"00",
		X"00",X"0C",X"B0",X"2D",X"81",X"00",X"00",X"05",X"C0",X"57",X"FF",X"FF",X"FF",X"FF",X"FD",X"FF",
		X"FA",X"00",X"AF",X"F2",X"6F",X"FF",X"D1",X"00",X"01",X"00",X"03",X"B0",X"F7",X"00",X"00",X"00",
		X"00",X"03",X"BC",X"FF",X"FF",X"FF",X"FF",X"FF",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"60",X"00",
		X"00",X"A0",X"03",X"0A",X"09",X"90",X"00",X"00",X"00",X"00",X"0F",X"FF",X"67",X"FF",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"C3",X"02",X"83",X"00",X"44",X"46",X"60",X"00",X"00",
		X"00",X"00",X"6F",X"F0",X"F0",X"54",X"79",X"7F",X"FF",X"DF",X"FF",X"FF",X"FF",X"FF",X"86",X"5B",
		X"FF",X"F0",X"3A",X"F4",X"BB",X"10",X"00",X"00",X"00",X"00",X"30",X"00",X"20",X"06",X"42",X"17",
		X"CB",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"4F",X"FF",X"F7",X"DF",X"FF",X"BE",X"30",X"00",X"22",
		X"20",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"4C",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",
		X"FA",X"79",X"FF",X"C0",X"00",X"00",X"04",X"87",X"C1",X"96",X"D0",X"03",X"00",X"00",X"00",X"00",
		X"2D",X"FF",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"43",X"00",X"00",X"00",X"06",
		X"20",X"AA",X"00",X"16",X"00",X"00",X"00",X"96",X"B0",X"40",X"07",X"FF",X"FF",X"6F",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"C6",X"00",X"03",X"88",X"90",X"00",X"00",X"00",X"00",X"6F",X"71",
		X"51",X"01",X"9D",X"F9",X"31",X"4F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A9",X"3E",X"FF",
		X"FF",X"A0",X"00",X"00",X"00",X"01",X"31",X"00",X"00",X"45",X"30",X"00",X"0E",X"FF",X"FF",X"FF",
		X"FF",X"FA",X"FF",X"FE",X"9C",X"BC",X"FF",X"FF",X"FC",X"10",X"24",X"10",X"01",X"07",X"00",X"01",
		X"00",X"00",X"00",X"00",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7E",
		X"30",X"08",X"60",X"00",X"59",X"C8",X"3B",X"D8",X"00",X"00",X"00",X"01",X"34",X"02",X"AF",X"AC",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"01",X"68",X"10",X"00",X"25",X"30",X"2B",X"60",
		X"00",X"00",X"37",X"93",X"50",X"3A",X"A5",X"27",X"32",X"6D",X"BC",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F7",X"37",X"A4",X"41",X"00",X"00",X"00",X"00",X"03",X"84",X"48",X"81",X"9E",X"C5",X"12",
		X"05",X"96",X"6F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"FF",X"FC",X"30",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"24",X"00",X"05",X"7E",X"CF",X"FF",X"FB",X"EF",X"FF",X"FE",X"BC",
		X"A8",X"8F",X"FF",X"FF",X"F9",X"87",X"63",X"27",X"78",X"50",X"00",X"30",X"00",X"00",X"00",X"00",
		X"5B",X"AF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CA",X"CF",X"FF",X"FF",X"C8",X"43",X"52",X"03",X"78",
		X"67",X"8A",X"CE",X"83",X"00",X"00",X"00",X"00",X"11",X"03",X"42",X"5B",X"FC",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"DB",X"BA",X"71",X"02",X"50",X"05",X"AB",X"87",X"00",X"00",X"03",X"73",X"13",
		X"67",X"10",X"01",X"10",X"00",X"45",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"B8",X"DD",X"74",
		X"9B",X"84",X"00",X"00",X"00",X"01",X"10",X"36",X"66",X"87",X"20",X"00",X"01",X"57",X"CF",X"FE",
		X"DE",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"A7",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"17",X"DF",X"FF",X"FF",X"FF",X"DF",X"FC",X"7A",X"CF",X"FF",X"FF",X"FF",
		X"EB",X"A9",X"67",X"AB",X"63",X"24",X"63",X"00",X"00",X"00",X"00",X"00",X"03",X"79",X"89",X"FF",
		X"FF",X"FF",X"FD",X"EF",X"FF",X"FF",X"FF",X"E6",X"34",X"55",X"78",X"77",X"6A",X"CE",X"EA",X"75",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"57",X"87",X"87",X"9F",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"C9",X"87",X"62",X"14",X"89",X"89",X"72",X"00",X"12",X"66",X"68",X"B9",X"30",X"01",X"00",X"00",
		X"00",X"03",X"9C",X"DF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A8",X"CF",X"D9",X"41",X"00",X"00",
		X"00",X"00",X"26",X"87",X"8A",X"86",X"32",X"00",X"13",X"6B",X"D8",X"57",X"BC",X"DF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FD",X"97",X"65",X"10",X"00",X"00",X"00",X"01",X"21",X"00",X"00",X"01",
		X"7B",X"CC",X"AA",X"CC",X"BC",X"CB",X"AB",X"CC",X"BE",X"FF",X"FF",X"FF",X"FE",X"DE",X"FF",X"96",
		X"67",X"87",X"66",X"43",X"00",X"00",X"00",X"00",X"12",X"23",X"7A",X"BA",X"BA",X"97",X"BF",X"FF",
		X"FF",X"FF",X"FD",X"CC",X"B9",X"9C",X"B8",X"7A",X"DD",X"CA",X"99",X"97",X"44",X"31",X"00",X"00",
		X"00",X"00",X"33",X"20",X"01",X"25",X"9D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"B9",X"66",X"79",
		X"BA",X"73",X"23",X"32",X"22",X"45",X"78",X"53",X"35",X"56",X"63",X"00",X"00",X"02",X"35",X"9C",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"83",X"10",X"00",X"00",X"02",X"42",X"13",
		X"45",X"66",X"63",X"11",X"34",X"64",X"33",X"78",X"77",X"9A",X"AC",X"ED",X"DD",X"EF",X"FF",X"FF",
		X"FF",X"FF",X"C9",X"63",X"32",X"33",X"20",X"01",X"10",X"00",X"00",X"03",X"56",X"76",X"79",X"AA",
		X"AA",X"A9",X"98",X"88",X"9A",X"BD",X"FF",X"FF",X"FF",X"FF",X"FC",X"BB",X"BB",X"BB",X"A9",X"86",
		X"30",X"00",X"00",X"01",X"00",X"01",X"35",X"78",X"89",X"89",X"BC",X"CD",X"FF",X"FF",X"FD",X"CC",
		X"DD",X"EC",X"86",X"79",X"9A",X"CE",X"ED",X"C9",X"75",X"31",X"13",X"31",X"00",X"11",X"20",X"00",
		X"00",X"03",X"68",X"AE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"AA",X"BB",X"97",X"78",X"88",X"76",
		X"55",X"44",X"56",X"55",X"68",X"88",X"62",X"00",X"00",X"00",X"01",X"36",X"8A",X"BB",X"CE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"DB",X"A9",X"54",X"33",X"10",X"11",X"23",X"68",X"98",X"64",X"34",
		X"43",X"33",X"34",X"56",X"67",X"76",X"67",X"87",X"68",X"BF",X"FF",X"FF",X"FF",X"FF",X"FE",X"CB",
		X"A9",X"76",X"42",X"23",X"32",X"10",X"00",X"02",X"12",X"33",X"68",X"99",X"9B",X"A9",X"99",X"86",
		X"47",X"AD",X"EE",X"DF",X"FF",X"ED",X"DD",X"DD",X"ED",X"DC",X"CB",X"B9",X"74",X"31",X"00",X"00",
		X"00",X"00",X"02",X"22",X"36",X"77",X"88",X"89",X"BD",X"FF",X"FF",X"FF",X"FF",X"DB",X"BA",X"9A",
		X"BC",X"EE",X"DE",X"DC",X"97",X"77",X"66",X"53",X"32",X"22",X"10",X"00",X"00",X"00",X"01",X"36",
		X"99",X"BC",X"EF",X"FF",X"FF",X"FF",X"DC",X"DC",X"DD",X"DD",X"CA",X"86",X"44",X"56",X"66",X"56",
		X"89",X"99",X"86",X"52",X"10",X"00",X"01",X"23",X"33",X"46",X"8A",X"BC",X"DE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"EC",X"A8",X"65",X"43",X"22",X"34",X"66",X"66",X"66",X"54",X"44",X"55",X"66",X"76",
		X"44",X"56",X"55",X"45",X"78",X"AB",X"DF",X"FF",X"FF",X"FF",X"FF",X"FE",X"CA",X"86",X"66",X"76",
		X"53",X"21",X"00",X"00",X"01",X"13",X"46",X"78",X"88",X"77",X"54",X"46",X"89",X"AB",X"BC",X"CD",
		X"DE",X"FF",X"EF",X"FF",X"ED",X"EE",X"FE",X"DB",X"98",X"65",X"42",X"10",X"00",X"00",X"12",X"34",
		X"44",X"43",X"24",X"57",X"9A",X"BC",X"DD",X"DC",X"CC",X"CC",X"BB",X"BC",X"BC",X"DD",X"DC",X"BB",
		X"BB",X"98",X"77",X"66",X"55",X"44",X"33",X"32",X"10",X"00",X"00",X"23",X"57",X"9B",X"DE",X"EE",
		X"EE",X"ED",X"ED",X"ED",X"EE",X"ED",X"B9",X"99",X"87",X"65",X"67",X"76",X"77",X"77",X"66",X"53",
		X"22",X"22",X"21",X"11",X"34",X"57",X"89",X"99",X"AB",X"CD",X"EF",X"FF",X"FF",X"FF",X"FE",X"CB",
		X"96",X"55",X"56",X"65",X"56",X"54",X"42",X"33",X"34",X"56",X"65",X"44",X"55",X"45",X"55",X"55",
		X"46",X"79",X"AC",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"CB",X"BB",X"98",X"76",X"52",X"00",X"00",
		X"11",X"23",X"43",X"56",X"76",X"65",X"56",X"66",X"67",X"88",X"89",X"AB",X"BC",X"DE",X"ED",X"CC",
		X"EF",X"FF",X"FF",X"ED",X"CB",X"97",X"43",X"32",X"11",X"12",X"33",X"44",X"32",X"23",X"46",X"66",
		X"89",X"AB",X"BC",X"CC",X"CC",X"BC",X"BA",X"AB",X"CC",X"CC",X"CC",X"CD",X"CB",X"A9",X"87",X"67",
		X"55",X"66",X"65",X"41",X"00",X"00",X"01",X"23",X"47",X"89",X"AB",X"CC",X"DC",X"CC",X"CD",X"DF",
		X"FF",X"ED",X"CC",X"CB",X"A8",X"99",X"66",X"77",X"78",X"89",X"87",X"65",X"43",X"11",X"11",X"12",
		X"33",X"35",X"54",X"66",X"77",X"9A",X"CE",X"FF",X"FF",X"FF",X"FF",X"FC",X"BB",X"A9",X"87",X"76",
		X"66",X"56",X"65",X"55",X"55",X"44",X"45",X"55",X"54",X"55",X"54",X"43",X"34",X"57",X"8A",X"BB",
		X"CE",X"FF",X"FE",X"EF",X"FF",X"FF",X"ED",X"BB",X"A9",X"65",X"43",X"33",X"33",X"32",X"33",X"45",
		X"56",X"77",X"65",X"55",X"56",X"66",X"78",X"89",X"BC",X"CC",X"CC",X"CB",X"CC",X"DE",X"FF",X"FF",
		X"DC",X"B9",X"77",X"66",X"43",X"33",X"33",X"32",X"11",X"11",X"23",X"34",X"56",X"88",X"9A",X"BC",
		X"CC",X"CB",X"BB",X"CC",X"CB",X"CD",X"DE",X"EE",X"DC",X"BB",X"A9",X"98",X"88",X"88",X"76",X"54",
		X"32",X"10",X"00",X"12",X"23",X"33",X"46",X"68",X"99",X"AA",X"BC",X"DE",X"FD",X"EF",X"FE",X"ED",
		X"CB",X"BA",X"98",X"77",X"89",X"AA",X"98",X"77",X"66",X"43",X"32",X"33",X"44",X"33",X"34",X"44",
		X"44",X"67",X"79",X"BC",X"DD",X"EF",X"FF",X"FF",X"FE",X"DC",X"AA",X"99",X"88",X"77",X"76",X"65",
		X"44",X"33",X"55",X"67",X"77",X"66",X"65",X"43",X"33",X"34",X"67",X"89",X"AB",X"CD",X"DD",X"DE",
		X"EF",X"EE",X"ED",X"DD",X"CB",X"A9",X"87",X"65",X"32",X"22",X"33",X"45",X"55",X"65",X"55",X"44",
		X"45",X"66",X"77",X"89",X"99",X"99",X"AA",X"AB",X"CC",X"DE",X"FF",X"FF",X"FE",X"DC",X"CA",X"97",
		X"65",X"55",X"44",X"33",X"33",X"33",X"22",X"12",X"34",X"56",X"67",X"89",X"99",X"99",X"99",X"9A",
		X"BB",X"CC",X"EF",X"ED",X"DD",X"DC",X"CB",X"AA",X"AA",X"A9",X"97",X"66",X"65",X"43",X"22",X"22",
		X"23",X"33",X"45",X"67",X"77",X"77",X"89",X"9A",X"BD",X"DE",X"EE",X"ED",X"CC",X"BA",X"99",X"99",
		X"AB",X"A9",X"98",X"77",X"65",X"44",X"34",X"44",X"44",X"44",X"44",X"44",X"44",X"45",X"67",X"89",
		X"AC",X"DE",X"EE",X"FF",X"EE",X"DC",X"CC",X"CC",X"CB",X"A9",X"87",X"65",X"44",X"44",X"45",X"55",
		X"66",X"65",X"54",X"43",X"44",X"45",X"56",X"67",X"89",X"9A",X"BC",X"CD",X"CD",X"DD",X"EF",X"FF",
		X"FF",X"EC",X"BA",X"86",X"54",X"44",X"44",X"44",X"55",X"54",X"43",X"34",X"44",X"55",X"66",X"77",
		X"77",X"78",X"89",X"99",X"AB",X"CC",X"DE",X"EF",X"FF",X"FE",X"DC",X"BA",X"99",X"88",X"77",X"66",
		X"54",X"33",X"21",X"22",X"33",X"45",X"67",X"87",X"88",X"77",X"88",X"99",X"AB",X"AC",X"CC",X"CD",
		X"DD",X"DC",X"CB",X"BB",X"BB",X"BA",X"A9",X"98",X"76",X"54",X"32",X"21",X"12",X"33",X"44",X"55",
		X"56",X"65",X"78",X"9A",X"BC",X"DD",X"DD",X"DD",X"DC",X"CC",X"BB",X"BB",X"BB",X"AA",X"AA",X"99",
		X"77",X"65",X"54",X"43",X"44",X"44",X"33",X"33",X"33",X"33",X"45",X"67",X"9A",X"AC",X"CD",X"DD",
		X"DD",X"DD",X"DD",X"DD",X"DC",X"CB",X"BA",X"98",X"77",X"66",X"66",X"66",X"66",X"66",X"54",X"44",
		X"33",X"33",X"34",X"56",X"68",X"89",X"99",X"9A",X"BB",X"CD",X"EE",X"FF",X"FF",X"ED",X"CB",X"A9",
		X"98",X"77",X"66",X"66",X"66",X"54",X"44",X"43",X"44",X"44",X"45",X"66",X"67",X"78",X"87",X"88",
		X"89",X"AB",X"CD",X"DE",X"EE",X"ED",X"DC",X"CB",X"BA",X"99",X"99",X"88",X"76",X"54",X"33",X"23",
		X"33",X"34",X"44",X"55",X"66",X"77",X"77",X"78",X"9A",X"AB",X"CC",X"DD",X"DD",X"DC",X"CC",X"CC",
		X"BB",X"BB",X"BB",X"B9",X"98",X"76",X"54",X"33",X"34",X"44",X"43",X"33",X"33",X"33",X"45",X"57",
		X"89",X"9A",X"BC",X"DD",X"DC",X"CC",X"CC",X"CB",X"CC",X"CC",X"CC",X"BA",X"A9",X"88",X"76",X"66",
		X"66",X"66",X"65",X"44",X"32",X"22",X"23",X"44",X"56",X"78",X"99",X"AB",X"BB",X"CC",X"CD",X"CD",
		X"DD",X"DD",X"DC",X"BA",X"99",X"77",X"76",X"77",X"77",X"77",X"76",X"65",X"44",X"33",X"34",X"45",
		X"56",X"66",X"77",X"77",X"89",X"AB",X"CC",X"DE",X"EF",X"EE",X"ED",X"CC",X"B9",X"98",X"88",X"87",
		X"76",X"66",X"55",X"44",X"44",X"44",X"44",X"55",X"66",X"66",X"65",X"56",X"67",X"89",X"9B",X"BC",
		X"DE",X"EE",X"EE",X"ED",X"CC",X"CB",X"BB",X"AA",X"98",X"77",X"65",X"43",X"33",X"34",X"43",X"44",
		X"55",X"54",X"55",X"56",X"66",X"78",X"89",X"AB",X"BB",X"CB",X"CC",X"CC",X"CC",X"DD",X"DD",X"DC",
		X"CB",X"99",X"77",X"66",X"55",X"55",X"44",X"43",X"44",X"43",X"33",X"44",X"55",X"67",X"89",X"99",
		X"AA",X"BB",X"BB",X"BB",X"CC",X"CD",X"DD",X"DC",X"CB",X"A9",X"88",X"78",X"87",X"76",X"70",X"70",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"70",X"70");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
